magic
tech sky130A
magscale 1 2
timestamp 1678386439
<< metal1 >>
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 397546 700312 397552 700324
rect 332560 700284 397552 700312
rect 332560 700272 332566 700284
rect 397546 700272 397552 700284
rect 397604 700272 397610 700324
rect 194686 700000 194692 700052
rect 194744 700040 194750 700052
rect 202782 700040 202788 700052
rect 194744 700012 202788 700040
rect 194744 700000 194750 700012
rect 202782 700000 202788 700012
rect 202840 700000 202846 700052
rect 260098 699660 260104 699712
rect 260156 699700 260162 699712
rect 267642 699700 267648 699712
rect 260156 699672 267648 699700
rect 260156 699660 260162 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 193122 696940 193128 696992
rect 193180 696980 193186 696992
rect 194686 696980 194692 696992
rect 193180 696952 194692 696980
rect 193180 696940 193186 696952
rect 194686 696940 194692 696952
rect 194744 696940 194750 696992
rect 188338 694152 188344 694204
rect 188396 694192 188402 694204
rect 193122 694192 193128 694204
rect 188396 694164 193128 694192
rect 188396 694152 188402 694164
rect 193122 694152 193128 694164
rect 193180 694152 193186 694204
rect 253934 690276 253940 690328
rect 253992 690316 253998 690328
rect 260098 690316 260104 690328
rect 253992 690288 260104 690316
rect 253992 690276 253998 690288
rect 260098 690276 260104 690288
rect 260156 690276 260162 690328
rect 238754 683748 238760 683800
rect 238812 683788 238818 683800
rect 253934 683788 253940 683800
rect 238812 683760 253940 683788
rect 238812 683748 238818 683760
rect 253934 683748 253940 683760
rect 253992 683748 253998 683800
rect 233878 679872 233884 679924
rect 233936 679912 233942 679924
rect 238754 679912 238760 679924
rect 233936 679884 238760 679912
rect 233936 679872 233942 679884
rect 238754 679872 238760 679884
rect 238812 679872 238818 679924
rect 183186 679056 183192 679108
rect 183244 679096 183250 679108
rect 188338 679096 188344 679108
rect 183244 679068 188344 679096
rect 183244 679056 183250 679068
rect 188338 679056 188344 679068
rect 188396 679056 188402 679108
rect 180058 677152 180064 677204
rect 180116 677192 180122 677204
rect 183186 677192 183192 677204
rect 180116 677164 183192 677192
rect 180116 677152 180122 677164
rect 183186 677152 183192 677164
rect 183244 677152 183250 677204
rect 175918 657160 175924 657212
rect 175976 657200 175982 657212
rect 180058 657200 180064 657212
rect 175976 657172 180064 657200
rect 175976 657160 175982 657172
rect 180058 657160 180064 657172
rect 180116 657160 180122 657212
rect 156598 643696 156604 643748
rect 156656 643736 156662 643748
rect 175918 643736 175924 643748
rect 156656 643708 175924 643736
rect 156656 643696 156662 643708
rect 175918 643696 175924 643708
rect 175976 643696 175982 643748
rect 150434 635468 150440 635520
rect 150492 635508 150498 635520
rect 156598 635508 156604 635520
rect 150492 635480 156604 635508
rect 150492 635468 150498 635480
rect 156598 635468 156604 635480
rect 156656 635468 156662 635520
rect 141418 631320 141424 631372
rect 141476 631360 141482 631372
rect 150434 631360 150440 631372
rect 141476 631332 150440 631360
rect 141476 631320 141482 631332
rect 150434 631320 150440 631332
rect 150492 631320 150498 631372
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 43438 605860 43444 605872
rect 3292 605832 43444 605860
rect 3292 605820 3298 605832
rect 43438 605820 43444 605832
rect 43496 605820 43502 605872
rect 211798 591268 211804 591320
rect 211856 591308 211862 591320
rect 233878 591308 233884 591320
rect 211856 591280 233884 591308
rect 211856 591268 211862 591280
rect 233878 591268 233884 591280
rect 233936 591268 233942 591320
rect 422938 590656 422944 590708
rect 422996 590696 423002 590708
rect 579706 590696 579712 590708
rect 422996 590668 579712 590696
rect 422996 590656 423002 590668
rect 579706 590656 579712 590668
rect 579764 590656 579770 590708
rect 209038 580932 209044 580984
rect 209096 580972 209102 580984
rect 211798 580972 211804 580984
rect 209096 580944 211804 580972
rect 209096 580932 209102 580944
rect 211798 580932 211804 580944
rect 211856 580932 211862 580984
rect 134794 574064 134800 574116
rect 134852 574104 134858 574116
rect 141418 574104 141424 574116
rect 134852 574076 141424 574104
rect 134852 574064 134858 574076
rect 141418 574064 141424 574076
rect 141476 574064 141482 574116
rect 127618 570936 127624 570988
rect 127676 570976 127682 570988
rect 134794 570976 134800 570988
rect 127676 570948 134800 570976
rect 127676 570936 127682 570948
rect 134794 570936 134800 570948
rect 134852 570936 134858 570988
rect 195238 570596 195244 570648
rect 195296 570636 195302 570648
rect 209038 570636 209044 570648
rect 195296 570608 209044 570636
rect 195296 570596 195302 570608
rect 209038 570596 209044 570608
rect 209096 570596 209102 570648
rect 189718 567808 189724 567860
rect 189776 567848 189782 567860
rect 195238 567848 195244 567860
rect 189776 567820 195244 567848
rect 189776 567808 189782 567820
rect 195238 567808 195244 567820
rect 195296 567808 195302 567860
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 43530 553432 43536 553444
rect 3384 553404 43536 553432
rect 3384 553392 3390 553404
rect 43530 553392 43536 553404
rect 43588 553392 43594 553444
rect 124858 552644 124864 552696
rect 124916 552684 124922 552696
rect 127618 552684 127624 552696
rect 124916 552656 127624 552684
rect 124916 552644 124922 552656
rect 127618 552644 127624 552656
rect 127676 552644 127682 552696
rect 396718 536800 396724 536852
rect 396776 536840 396782 536852
rect 580166 536840 580172 536852
rect 396776 536812 580172 536840
rect 396776 536800 396782 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 119338 532040 119344 532092
rect 119396 532080 119402 532092
rect 124858 532080 124864 532092
rect 119396 532052 124864 532080
rect 119396 532040 119402 532052
rect 124858 532040 124864 532052
rect 124916 532040 124922 532092
rect 184382 511912 184388 511964
rect 184440 511952 184446 511964
rect 189718 511952 189724 511964
rect 184440 511924 189724 511952
rect 184440 511912 184446 511924
rect 189718 511912 189724 511924
rect 189776 511912 189782 511964
rect 114554 511164 114560 511216
rect 114612 511204 114618 511216
rect 119338 511204 119344 511216
rect 114612 511176 119344 511204
rect 114612 511164 114618 511176
rect 119338 511164 119344 511176
rect 119396 511164 119402 511216
rect 117958 508512 117964 508564
rect 118016 508552 118022 508564
rect 137830 508552 137836 508564
rect 118016 508524 137836 508552
rect 118016 508512 118022 508524
rect 137830 508512 137836 508524
rect 137888 508512 137894 508564
rect 178678 507084 178684 507136
rect 178736 507124 178742 507136
rect 184382 507124 184388 507136
rect 178736 507096 184388 507124
rect 178736 507084 178742 507096
rect 184382 507084 184388 507096
rect 184440 507084 184446 507136
rect 112438 504160 112444 504212
rect 112496 504200 112502 504212
rect 114554 504200 114560 504212
rect 112496 504172 114560 504200
rect 112496 504160 112502 504172
rect 114554 504160 114560 504172
rect 114612 504160 114618 504212
rect 116578 487160 116584 487212
rect 116636 487200 116642 487212
rect 117958 487200 117964 487212
rect 116636 487172 117964 487200
rect 116636 487160 116642 487172
rect 117958 487160 117964 487172
rect 118016 487160 118022 487212
rect 418798 484372 418804 484424
rect 418856 484412 418862 484424
rect 580166 484412 580172 484424
rect 418856 484384 580172 484412
rect 418856 484372 418862 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 174538 482944 174544 482996
rect 174596 482984 174602 482996
rect 178678 482984 178684 482996
rect 174596 482956 178684 482984
rect 174596 482944 174602 482956
rect 178678 482944 178684 482956
rect 178736 482944 178742 482996
rect 115198 472948 115204 473000
rect 115256 472988 115262 473000
rect 116578 472988 116584 473000
rect 115256 472960 116584 472988
rect 115256 472948 115262 472960
rect 116578 472948 116584 472960
rect 116636 472948 116642 473000
rect 166258 467100 166264 467152
rect 166316 467140 166322 467152
rect 174538 467140 174544 467152
rect 166316 467112 174544 467140
rect 166316 467100 166322 467112
rect 174538 467100 174544 467112
rect 174596 467100 174602 467152
rect 93118 461592 93124 461644
rect 93176 461632 93182 461644
rect 112438 461632 112444 461644
rect 93176 461604 112444 461632
rect 93176 461592 93182 461604
rect 112438 461592 112444 461604
rect 112496 461592 112502 461644
rect 162854 452820 162860 452872
rect 162912 452860 162918 452872
rect 166258 452860 166264 452872
rect 162912 452832 166264 452860
rect 162912 452820 162918 452832
rect 166258 452820 166264 452832
rect 166316 452820 166322 452872
rect 2774 449488 2780 449540
rect 2832 449528 2838 449540
rect 4890 449528 4896 449540
rect 2832 449500 4896 449528
rect 2832 449488 2838 449500
rect 4890 449488 4896 449500
rect 4948 449488 4954 449540
rect 155218 447040 155224 447092
rect 155276 447080 155282 447092
rect 162854 447080 162860 447092
rect 155276 447052 162860 447080
rect 155276 447040 155282 447052
rect 162854 447040 162860 447052
rect 162912 447040 162918 447092
rect 442258 444388 442264 444440
rect 442316 444428 442322 444440
rect 580166 444428 580172 444440
rect 442316 444400 580172 444428
rect 442316 444388 442322 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 79318 436704 79324 436756
rect 79376 436744 79382 436756
rect 93118 436744 93124 436756
rect 79376 436716 93124 436744
rect 79376 436704 79382 436716
rect 93118 436704 93124 436716
rect 93176 436704 93182 436756
rect 413278 430584 413284 430636
rect 413336 430624 413342 430636
rect 580166 430624 580172 430636
rect 413336 430596 580172 430624
rect 413336 430584 413342 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 76926 419500 76932 419552
rect 76984 419540 76990 419552
rect 79318 419540 79324 419552
rect 76984 419512 79324 419540
rect 76984 419500 76990 419512
rect 79318 419500 79324 419512
rect 79376 419500 79382 419552
rect 73154 417800 73160 417852
rect 73212 417840 73218 417852
rect 76926 417840 76932 417852
rect 73212 417812 76932 417840
rect 73212 417800 73218 417812
rect 76926 417800 76932 417812
rect 76984 417800 76990 417852
rect 64138 413244 64144 413296
rect 64196 413284 64202 413296
rect 73154 413284 73160 413296
rect 64196 413256 73160 413284
rect 64196 413244 64202 413256
rect 73154 413244 73160 413256
rect 73212 413244 73218 413296
rect 152458 411272 152464 411324
rect 152516 411312 152522 411324
rect 155218 411312 155224 411324
rect 152516 411284 155224 411312
rect 152516 411272 152522 411284
rect 155218 411272 155224 411284
rect 155276 411272 155282 411324
rect 50982 404948 50988 405000
rect 51040 404988 51046 405000
rect 64138 404988 64144 405000
rect 51040 404960 64144 404988
rect 51040 404948 51046 404960
rect 64138 404948 64144 404960
rect 64196 404948 64202 405000
rect 47578 401616 47584 401668
rect 47636 401656 47642 401668
rect 50982 401656 50988 401668
rect 47636 401628 50988 401656
rect 47636 401616 47642 401628
rect 50982 401616 50988 401628
rect 51040 401616 51046 401668
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 13078 397508 13084 397520
rect 3384 397480 13084 397508
rect 3384 397468 3390 397480
rect 13078 397468 13084 397480
rect 13136 397468 13142 397520
rect 46198 382236 46204 382288
rect 46256 382276 46262 382288
rect 47578 382276 47584 382288
rect 46256 382248 47584 382276
rect 46256 382236 46262 382248
rect 47578 382236 47584 382248
rect 47636 382236 47642 382288
rect 421558 378156 421564 378208
rect 421616 378196 421622 378208
rect 580166 378196 580172 378208
rect 421616 378168 580172 378196
rect 421616 378156 421622 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 115290 363604 115296 363656
rect 115348 363644 115354 363656
rect 152458 363644 152464 363656
rect 115348 363616 152464 363644
rect 115348 363604 115354 363616
rect 152458 363604 152464 363616
rect 152516 363604 152522 363656
rect 58618 356668 58624 356720
rect 58676 356708 58682 356720
rect 115198 356708 115204 356720
rect 58676 356680 115204 356708
rect 58676 356668 58682 356680
rect 115198 356668 115204 356680
rect 115256 356668 115262 356720
rect 45186 350072 45192 350124
rect 45244 350112 45250 350124
rect 46198 350112 46204 350124
rect 45244 350084 46204 350112
rect 45244 350072 45250 350084
rect 46198 350072 46204 350084
rect 46256 350072 46262 350124
rect 2774 345176 2780 345228
rect 2832 345216 2838 345228
rect 5074 345216 5080 345228
rect 2832 345188 5080 345216
rect 2832 345176 2838 345188
rect 5074 345176 5080 345188
rect 5132 345176 5138 345228
rect 57238 339668 57244 339720
rect 57296 339708 57302 339720
rect 58618 339708 58624 339720
rect 57296 339680 58624 339708
rect 57296 339668 57302 339680
rect 58618 339668 58624 339680
rect 58676 339668 58682 339720
rect 95234 337356 95240 337408
rect 95292 337396 95298 337408
rect 115290 337396 115296 337408
rect 95292 337368 115296 337396
rect 95292 337356 95298 337368
rect 115290 337356 115296 337368
rect 115348 337356 115354 337408
rect 93118 328856 93124 328908
rect 93176 328896 93182 328908
rect 95234 328896 95240 328908
rect 93176 328868 95240 328896
rect 93176 328856 93182 328868
rect 95234 328856 95240 328868
rect 95292 328856 95298 328908
rect 55950 327020 55956 327072
rect 56008 327060 56014 327072
rect 57238 327060 57244 327072
rect 56008 327032 57244 327060
rect 56008 327020 56014 327032
rect 57238 327020 57244 327032
rect 57296 327020 57302 327072
rect 417418 324300 417424 324352
rect 417476 324340 417482 324352
rect 579614 324340 579620 324352
rect 417476 324312 579620 324340
rect 417476 324300 417482 324312
rect 579614 324300 579620 324312
rect 579672 324300 579678 324352
rect 54478 321104 54484 321156
rect 54536 321144 54542 321156
rect 55950 321144 55956 321156
rect 54536 321116 55956 321144
rect 54536 321104 54542 321116
rect 55950 321104 55956 321116
rect 56008 321104 56014 321156
rect 53098 309068 53104 309120
rect 53156 309108 53162 309120
rect 54478 309108 54484 309120
rect 53156 309080 54484 309108
rect 53156 309068 53162 309080
rect 54478 309068 54484 309080
rect 54536 309068 54542 309120
rect 87598 304988 87604 305040
rect 87656 305028 87662 305040
rect 93118 305028 93124 305040
rect 87656 305000 93124 305028
rect 87656 304988 87662 305000
rect 93118 304988 93124 305000
rect 93176 304988 93182 305040
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 43622 292584 43628 292596
rect 3384 292556 43628 292584
rect 3384 292544 3390 292556
rect 43622 292544 43628 292556
rect 43680 292544 43686 292596
rect 73154 287648 73160 287700
rect 73212 287688 73218 287700
rect 87598 287688 87604 287700
rect 73212 287660 87604 287688
rect 73212 287648 73218 287660
rect 87598 287648 87604 287660
rect 87656 287648 87662 287700
rect 57882 280780 57888 280832
rect 57940 280820 57946 280832
rect 73154 280820 73160 280832
rect 57940 280792 73160 280820
rect 57940 280780 57946 280792
rect 73154 280780 73160 280792
rect 73212 280780 73218 280832
rect 51074 279420 51080 279472
rect 51132 279460 51138 279472
rect 53098 279460 53104 279472
rect 51132 279432 53104 279460
rect 51132 279420 51138 279432
rect 53098 279420 53104 279432
rect 53156 279420 53162 279472
rect 47578 277992 47584 278044
rect 47636 278032 47642 278044
rect 57882 278032 57888 278044
rect 47636 278004 57888 278032
rect 47636 277992 47642 278004
rect 57882 277992 57888 278004
rect 57940 277992 57946 278044
rect 48958 273232 48964 273284
rect 49016 273272 49022 273284
rect 50982 273272 50988 273284
rect 49016 273244 50988 273272
rect 49016 273232 49022 273244
rect 50982 273232 50988 273244
rect 51040 273232 51046 273284
rect 410518 271872 410524 271924
rect 410576 271912 410582 271924
rect 579614 271912 579620 271924
rect 410576 271884 579620 271912
rect 410576 271872 410582 271884
rect 579614 271872 579620 271884
rect 579672 271872 579678 271924
rect 46198 270172 46204 270224
rect 46256 270212 46262 270224
rect 47578 270212 47584 270224
rect 46256 270184 47584 270212
rect 46256 270172 46262 270184
rect 47578 270172 47584 270184
rect 47636 270172 47642 270224
rect 47670 262216 47676 262268
rect 47728 262256 47734 262268
rect 48958 262256 48964 262268
rect 47728 262228 48964 262256
rect 47728 262216 47734 262228
rect 48958 262216 48964 262228
rect 49016 262216 49022 262268
rect 46290 259224 46296 259276
rect 46348 259264 46354 259276
rect 47670 259264 47676 259276
rect 46348 259236 47676 259264
rect 46348 259224 46354 259236
rect 47670 259224 47676 259236
rect 47728 259224 47734 259276
rect 45278 249772 45284 249824
rect 45336 249812 45342 249824
rect 46290 249812 46296 249824
rect 45336 249784 46296 249812
rect 45336 249772 45342 249784
rect 46290 249772 46296 249784
rect 46348 249772 46354 249824
rect 3326 240116 3332 240168
rect 3384 240156 3390 240168
rect 21358 240156 21364 240168
rect 3384 240128 21364 240156
rect 3384 240116 3390 240128
rect 21358 240116 21364 240128
rect 21416 240116 21422 240168
rect 44818 225972 44824 226024
rect 44876 226012 44882 226024
rect 72970 226012 72976 226024
rect 44876 225984 72976 226012
rect 44876 225972 44882 225984
rect 72970 225972 72976 225984
rect 73028 225972 73034 226024
rect 45002 224952 45008 225004
rect 45060 224992 45066 225004
rect 68922 224992 68928 225004
rect 45060 224964 68928 224992
rect 45060 224952 45066 224964
rect 68922 224952 68928 224964
rect 68980 224952 68986 225004
rect 45462 224000 45468 224052
rect 45520 224040 45526 224052
rect 46198 224040 46204 224052
rect 45520 224012 46204 224040
rect 45520 224000 45526 224012
rect 46198 224000 46204 224012
rect 46256 224000 46262 224052
rect 45278 215908 45284 215960
rect 45336 215948 45342 215960
rect 56686 215948 56692 215960
rect 45336 215920 56692 215948
rect 45336 215908 45342 215920
rect 56686 215908 56692 215920
rect 56744 215908 56750 215960
rect 57330 215908 57336 215960
rect 57388 215948 57394 215960
rect 68278 215948 68284 215960
rect 57388 215920 68284 215948
rect 57388 215908 57394 215920
rect 68278 215908 68284 215920
rect 68336 215908 68342 215960
rect 45186 214548 45192 214600
rect 45244 214588 45250 214600
rect 45244 214560 45554 214588
rect 45244 214548 45250 214560
rect 45526 214316 45554 214560
rect 57790 214316 57796 214328
rect 45526 214288 57796 214316
rect 57790 214276 57796 214288
rect 57848 214276 57854 214328
rect 174538 211080 174544 211132
rect 174596 211120 174602 211132
rect 176654 211120 176660 211132
rect 174596 211092 176660 211120
rect 174596 211080 174602 211092
rect 176654 211080 176660 211092
rect 176712 211080 176718 211132
rect 177298 210400 177304 210452
rect 177356 210440 177362 210452
rect 580350 210440 580356 210452
rect 177356 210412 580356 210440
rect 177356 210400 177362 210412
rect 580350 210400 580356 210412
rect 580408 210400 580414 210452
rect 45462 209924 45468 209976
rect 45520 209964 45526 209976
rect 47578 209964 47584 209976
rect 45520 209936 47584 209964
rect 45520 209924 45526 209936
rect 47578 209924 47584 209936
rect 47636 209924 47642 209976
rect 57790 209040 57796 209092
rect 57848 209080 57854 209092
rect 69658 209080 69664 209092
rect 57848 209052 69664 209080
rect 57848 209040 57854 209052
rect 69658 209040 69664 209052
rect 69716 209040 69722 209092
rect 68278 208904 68284 208956
rect 68336 208944 68342 208956
rect 75546 208944 75552 208956
rect 68336 208916 75552 208944
rect 68336 208904 68342 208916
rect 75546 208904 75552 208916
rect 75604 208904 75610 208956
rect 69658 204892 69664 204944
rect 69716 204932 69722 204944
rect 85114 204932 85120 204944
rect 69716 204904 85120 204932
rect 69716 204892 69722 204904
rect 85114 204892 85120 204904
rect 85172 204892 85178 204944
rect 47578 202784 47584 202836
rect 47636 202824 47642 202836
rect 51718 202824 51724 202836
rect 47636 202796 51724 202824
rect 47636 202784 47642 202796
rect 51718 202784 51724 202796
rect 51776 202784 51782 202836
rect 75546 201492 75552 201544
rect 75604 201532 75610 201544
rect 75604 201504 75960 201532
rect 75604 201492 75610 201504
rect 75932 201464 75960 201504
rect 78030 201464 78036 201476
rect 75932 201436 78036 201464
rect 78030 201424 78036 201436
rect 78088 201424 78094 201476
rect 85114 201424 85120 201476
rect 85172 201464 85178 201476
rect 87598 201464 87604 201476
rect 85172 201436 87604 201464
rect 85172 201424 85178 201436
rect 87598 201424 87604 201436
rect 87656 201424 87662 201476
rect 78030 198704 78036 198756
rect 78088 198744 78094 198756
rect 78088 198716 80100 198744
rect 78088 198704 78094 198716
rect 80072 198676 80100 198716
rect 81434 198676 81440 198688
rect 80072 198648 81440 198676
rect 81434 198636 81440 198648
rect 81492 198636 81498 198688
rect 81434 194556 81440 194608
rect 81492 194596 81498 194608
rect 81492 194568 84194 194596
rect 81492 194556 81498 194568
rect 84166 194528 84194 194568
rect 84838 194528 84844 194540
rect 84166 194500 84844 194528
rect 84838 194488 84844 194500
rect 84896 194488 84902 194540
rect 87598 194488 87604 194540
rect 87656 194528 87662 194540
rect 89714 194528 89720 194540
rect 87656 194500 89720 194528
rect 87656 194488 87662 194500
rect 89714 194488 89720 194500
rect 89772 194488 89778 194540
rect 89714 191088 89720 191140
rect 89772 191128 89778 191140
rect 111058 191128 111064 191140
rect 89772 191100 111064 191128
rect 89772 191088 89778 191100
rect 111058 191088 111064 191100
rect 111116 191088 111122 191140
rect 149514 191088 149520 191140
rect 149572 191128 149578 191140
rect 266354 191128 266360 191140
rect 149572 191100 266360 191128
rect 149572 191088 149578 191100
rect 266354 191088 266360 191100
rect 266412 191088 266418 191140
rect 147582 189728 147588 189780
rect 147640 189768 147646 189780
rect 235994 189768 236000 189780
rect 147640 189740 236000 189768
rect 147640 189728 147646 189740
rect 235994 189728 236000 189740
rect 236052 189728 236058 189780
rect 146202 188300 146208 188352
rect 146260 188340 146266 188352
rect 207014 188340 207020 188352
rect 146260 188312 207020 188340
rect 146260 188300 146266 188312
rect 207014 188300 207020 188312
rect 207072 188300 207078 188352
rect 3142 187688 3148 187740
rect 3200 187728 3206 187740
rect 112438 187728 112444 187740
rect 3200 187700 112444 187728
rect 3200 187688 3206 187700
rect 112438 187688 112444 187700
rect 112496 187688 112502 187740
rect 144730 185580 144736 185632
rect 144788 185620 144794 185632
rect 174538 185620 174544 185632
rect 144788 185592 174544 185620
rect 144788 185580 144794 185592
rect 174538 185580 174544 185592
rect 174596 185580 174602 185632
rect 84838 184832 84844 184884
rect 84896 184872 84902 184884
rect 86218 184872 86224 184884
rect 84896 184844 86224 184872
rect 84896 184832 84902 184844
rect 86218 184832 86224 184844
rect 86276 184832 86282 184884
rect 134518 183948 134524 184000
rect 134576 183988 134582 184000
rect 137278 183988 137284 184000
rect 134576 183960 137284 183988
rect 134576 183948 134582 183960
rect 137278 183948 137284 183960
rect 137336 183948 137342 184000
rect 111058 182724 111064 182776
rect 111116 182764 111122 182776
rect 113542 182764 113548 182776
rect 111116 182736 113548 182764
rect 111116 182724 111122 182736
rect 113542 182724 113548 182736
rect 113600 182724 113606 182776
rect 151538 182452 151544 182504
rect 151596 182492 151602 182504
rect 154482 182492 154488 182504
rect 151596 182464 154488 182492
rect 151596 182452 151602 182464
rect 154482 182452 154488 182464
rect 154540 182452 154546 182504
rect 138566 182384 138572 182436
rect 138624 182424 138630 182436
rect 154666 182424 154672 182436
rect 138624 182396 154672 182424
rect 138624 182384 138630 182396
rect 154666 182384 154672 182396
rect 154724 182384 154730 182436
rect 133230 181976 133236 182028
rect 133288 182016 133294 182028
rect 136634 182016 136640 182028
rect 133288 181988 136640 182016
rect 133288 181976 133294 181988
rect 136634 181976 136640 181988
rect 136692 181976 136698 182028
rect 146018 181568 146024 181620
rect 146076 181568 146082 181620
rect 136542 181500 136548 181552
rect 136600 181540 136606 181552
rect 136600 181512 138322 181540
rect 136600 181500 136606 181512
rect 138216 181376 138414 181404
rect 118602 181160 118608 181212
rect 118660 181200 118666 181212
rect 138014 181200 138020 181212
rect 118660 181172 138020 181200
rect 118660 181160 118666 181172
rect 138014 181160 138020 181172
rect 138072 181160 138078 181212
rect 113818 181092 113824 181144
rect 113876 181132 113882 181144
rect 137830 181132 137836 181144
rect 113876 181104 137836 181132
rect 113876 181092 113882 181104
rect 137830 181092 137836 181104
rect 137888 181092 137894 181144
rect 137922 181092 137928 181144
rect 137980 181132 137986 181144
rect 138216 181132 138244 181376
rect 137980 181104 138244 181132
rect 137980 181092 137986 181104
rect 138014 181024 138020 181076
rect 138072 181064 138078 181076
rect 138492 181064 138520 181322
rect 138072 181036 138520 181064
rect 138072 181024 138078 181036
rect 128262 180956 128268 181008
rect 128320 180996 128326 181008
rect 128320 180968 138060 180996
rect 128320 180956 128326 180968
rect 138032 180928 138060 180968
rect 138860 180928 138888 181050
rect 138032 180900 138888 180928
rect 146018 180820 146024 180872
rect 146076 180820 146082 180872
rect 113542 180684 113548 180736
rect 113600 180724 113606 180736
rect 116578 180724 116584 180736
rect 113600 180696 116584 180724
rect 113600 180684 113606 180696
rect 116578 180684 116584 180696
rect 116636 180684 116642 180736
rect 146036 180600 146064 180820
rect 146018 180548 146024 180600
rect 146076 180548 146082 180600
rect 155494 180480 155500 180532
rect 155552 180520 155558 180532
rect 161474 180520 161480 180532
rect 155552 180492 161480 180520
rect 155552 180480 155558 180492
rect 161474 180480 161480 180492
rect 161532 180480 161538 180532
rect 155770 180412 155776 180464
rect 155828 180452 155834 180464
rect 163498 180452 163504 180464
rect 155828 180424 163504 180452
rect 155828 180412 155834 180424
rect 163498 180412 163504 180424
rect 163556 180412 163562 180464
rect 155402 180344 155408 180396
rect 155460 180384 155466 180396
rect 163590 180384 163596 180396
rect 155460 180356 163596 180384
rect 155460 180344 155466 180356
rect 163590 180344 163596 180356
rect 163648 180344 163654 180396
rect 129642 179460 129648 179512
rect 129700 179500 129706 179512
rect 136358 179500 136364 179512
rect 129700 179472 136364 179500
rect 129700 179460 129706 179472
rect 136358 179460 136364 179472
rect 136416 179460 136422 179512
rect 86218 179392 86224 179444
rect 86276 179432 86282 179444
rect 86276 179404 87000 179432
rect 86276 179392 86282 179404
rect 86972 179364 87000 179404
rect 133230 179392 133236 179444
rect 133288 179432 133294 179444
rect 140958 179432 140964 179444
rect 133288 179404 140964 179432
rect 133288 179392 133294 179404
rect 140958 179392 140964 179404
rect 141016 179392 141022 179444
rect 89438 179364 89444 179376
rect 86972 179336 89444 179364
rect 89438 179324 89444 179336
rect 89496 179324 89502 179376
rect 120718 178644 120724 178696
rect 120776 178684 120782 178696
rect 136542 178684 136548 178696
rect 120776 178656 136548 178684
rect 120776 178644 120782 178656
rect 136542 178644 136548 178656
rect 136600 178644 136606 178696
rect 162762 177828 162768 177880
rect 162820 177868 162826 177880
rect 164878 177868 164884 177880
rect 162820 177840 164884 177868
rect 162820 177828 162826 177840
rect 164878 177828 164884 177840
rect 164936 177828 164942 177880
rect 154666 177800 154672 177812
rect 154592 177772 154672 177800
rect 154592 177528 154620 177772
rect 154666 177760 154672 177772
rect 154724 177760 154730 177812
rect 154592 177500 154896 177528
rect 121362 177284 121368 177336
rect 121420 177324 121426 177336
rect 137922 177324 137928 177336
rect 121420 177296 137928 177324
rect 121420 177284 121426 177296
rect 137922 177284 137928 177296
rect 137980 177284 137986 177336
rect 154868 177324 154896 177500
rect 154868 177296 154988 177324
rect 141510 177012 141516 177064
rect 141568 177052 141574 177064
rect 146294 177052 146300 177064
rect 141568 177024 146300 177052
rect 141568 177012 141574 177024
rect 146294 177012 146300 177024
rect 146352 177012 146358 177064
rect 154960 176970 154988 177296
rect 161474 176468 161480 176520
rect 161532 176468 161538 176520
rect 161492 175908 161520 176468
rect 124858 175856 124864 175908
rect 124916 175896 124922 175908
rect 138566 175896 138572 175908
rect 124916 175868 138572 175896
rect 124916 175856 124922 175868
rect 138566 175856 138572 175868
rect 138624 175856 138630 175908
rect 161474 175856 161480 175908
rect 161532 175856 161538 175908
rect 161382 174972 161388 175024
rect 161440 174972 161446 175024
rect 161400 174752 161428 174972
rect 161382 174700 161388 174752
rect 161440 174700 161446 174752
rect 89438 173816 89444 173868
rect 89496 173856 89502 173868
rect 92474 173856 92480 173868
rect 89496 173828 92480 173856
rect 89496 173816 89502 173828
rect 92474 173816 92480 173828
rect 92532 173816 92538 173868
rect 161474 167560 161480 167612
rect 161532 167560 161538 167612
rect 161492 167340 161520 167560
rect 161474 167288 161480 167340
rect 161532 167288 161538 167340
rect 92474 167016 92480 167068
rect 92532 167056 92538 167068
rect 92532 167028 93854 167056
rect 92532 167016 92538 167028
rect 93826 166988 93854 167028
rect 95878 166988 95884 167000
rect 93826 166960 95884 166988
rect 95878 166948 95884 166960
rect 95936 166948 95942 167000
rect 51718 164840 51724 164892
rect 51776 164880 51782 164892
rect 66898 164880 66904 164892
rect 51776 164852 66904 164880
rect 51776 164840 51782 164852
rect 66898 164840 66904 164852
rect 66956 164840 66962 164892
rect 147490 162596 147496 162648
rect 147548 162596 147554 162648
rect 136450 161440 136456 161492
rect 136508 161480 136514 161492
rect 137830 161480 137836 161492
rect 136508 161452 137836 161480
rect 136508 161440 136514 161452
rect 137830 161440 137836 161452
rect 137888 161440 137894 161492
rect 147508 161276 147536 162596
rect 161474 161712 161480 161764
rect 161532 161712 161538 161764
rect 161492 161492 161520 161712
rect 163222 161576 163228 161628
rect 163280 161616 163286 161628
rect 164234 161616 164240 161628
rect 163280 161588 164240 161616
rect 163280 161576 163286 161588
rect 164234 161576 164240 161588
rect 164292 161576 164298 161628
rect 160462 161480 160468 161492
rect 151556 161452 160468 161480
rect 151556 161276 151584 161452
rect 160462 161440 160468 161452
rect 160520 161440 160526 161492
rect 161474 161440 161480 161492
rect 161532 161440 161538 161492
rect 147508 161248 151584 161276
rect 135438 161168 135444 161220
rect 135496 161208 135502 161220
rect 136450 161208 136456 161220
rect 135496 161180 136456 161208
rect 135496 161168 135502 161180
rect 136450 161168 136456 161180
rect 136508 161168 136514 161220
rect 163314 159332 163320 159384
rect 163372 159372 163378 159384
rect 173894 159372 173900 159384
rect 163372 159344 173900 159372
rect 163372 159332 163378 159344
rect 173894 159332 173900 159344
rect 173952 159332 173958 159384
rect 133782 158720 133788 158772
rect 133840 158760 133846 158772
rect 136634 158760 136640 158772
rect 133840 158732 136640 158760
rect 133840 158720 133846 158732
rect 136634 158720 136640 158732
rect 136692 158720 136698 158772
rect 132402 158040 132408 158092
rect 132460 158080 132466 158092
rect 135622 158080 135628 158092
rect 132460 158052 135628 158080
rect 132460 158040 132466 158052
rect 135622 158040 135628 158052
rect 135680 158040 135686 158092
rect 131022 157360 131028 157412
rect 131080 157400 131086 157412
rect 134518 157400 134524 157412
rect 131080 157372 134524 157400
rect 131080 157360 131086 157372
rect 134518 157360 134524 157372
rect 134576 157360 134582 157412
rect 136542 157360 136548 157412
rect 136600 157400 136606 157412
rect 138658 157400 138664 157412
rect 136600 157372 138664 157400
rect 136600 157360 136606 157372
rect 138658 157360 138664 157372
rect 138716 157360 138722 157412
rect 151354 157360 151360 157412
rect 151412 157400 151418 157412
rect 152458 157400 152464 157412
rect 151412 157372 152464 157400
rect 151412 157360 151418 157372
rect 152458 157360 152464 157372
rect 152516 157360 152522 157412
rect 66898 155864 66904 155916
rect 66956 155904 66962 155916
rect 69290 155904 69296 155916
rect 66956 155876 69296 155904
rect 66956 155864 66962 155876
rect 69290 155864 69296 155876
rect 69348 155864 69354 155916
rect 95878 155864 95884 155916
rect 95936 155904 95942 155916
rect 97258 155904 97264 155916
rect 95936 155876 97264 155904
rect 95936 155864 95942 155876
rect 97258 155864 97264 155876
rect 97316 155864 97322 155916
rect 148502 155728 148508 155780
rect 148560 155768 148566 155780
rect 148962 155768 148968 155780
rect 148560 155740 148968 155768
rect 148560 155728 148566 155740
rect 148962 155728 148968 155740
rect 149020 155728 149026 155780
rect 69290 152464 69296 152516
rect 69348 152504 69354 152516
rect 84194 152504 84200 152516
rect 69348 152476 84200 152504
rect 69348 152464 69354 152476
rect 84194 152464 84200 152476
rect 84252 152464 84258 152516
rect 84194 149064 84200 149116
rect 84252 149104 84258 149116
rect 87598 149104 87604 149116
rect 84252 149076 87604 149104
rect 84252 149064 84258 149076
rect 87598 149064 87604 149076
rect 87656 149064 87662 149116
rect 164878 146208 164884 146260
rect 164936 146248 164942 146260
rect 165890 146248 165896 146260
rect 164936 146220 165896 146248
rect 164936 146208 164942 146220
rect 165890 146208 165896 146220
rect 165948 146208 165954 146260
rect 124030 137912 124036 137964
rect 124088 137952 124094 137964
rect 124858 137952 124864 137964
rect 124088 137924 124864 137952
rect 124088 137912 124094 137924
rect 124858 137912 124864 137924
rect 124916 137912 124922 137964
rect 146202 137912 146208 137964
rect 146260 137952 146266 137964
rect 147490 137952 147496 137964
rect 146260 137924 147496 137952
rect 146260 137912 146266 137924
rect 147490 137912 147496 137924
rect 147548 137912 147554 137964
rect 152458 137912 152464 137964
rect 152516 137952 152522 137964
rect 155310 137952 155316 137964
rect 152516 137924 155316 137952
rect 152516 137912 152522 137924
rect 155310 137912 155316 137924
rect 155368 137912 155374 137964
rect 134978 137844 134984 137896
rect 135036 137884 135042 137896
rect 136450 137884 136456 137896
rect 135036 137856 136456 137884
rect 135036 137844 135042 137856
rect 136450 137844 136456 137856
rect 136508 137844 136514 137896
rect 150342 137844 150348 137896
rect 150400 137884 150406 137896
rect 153746 137884 153752 137896
rect 150400 137856 153752 137884
rect 150400 137844 150406 137856
rect 153746 137844 153752 137856
rect 153804 137844 153810 137896
rect 148870 137776 148876 137828
rect 148928 137816 148934 137828
rect 152182 137816 152188 137828
rect 148928 137788 152188 137816
rect 148928 137776 148934 137788
rect 152182 137776 152188 137788
rect 152240 137776 152246 137828
rect 156874 137640 156880 137692
rect 156932 137680 156938 137692
rect 163590 137680 163596 137692
rect 156932 137652 163596 137680
rect 156932 137640 156938 137652
rect 163590 137640 163596 137652
rect 163648 137640 163654 137692
rect 161382 137300 161388 137352
rect 161440 137340 161446 137352
rect 170950 137340 170956 137352
rect 161440 137312 170956 137340
rect 161440 137300 161446 137312
rect 170950 137300 170956 137312
rect 171008 137300 171014 137352
rect 162762 137232 162768 137284
rect 162820 137272 162826 137284
rect 172514 137272 172520 137284
rect 162820 137244 172520 137272
rect 162820 137232 162826 137244
rect 172514 137232 172520 137244
rect 172572 137232 172578 137284
rect 158438 137096 158444 137148
rect 158496 137136 158502 137148
rect 163498 137136 163504 137148
rect 158496 137108 163504 137136
rect 158496 137096 158502 137108
rect 163498 137096 163504 137108
rect 163556 137096 163562 137148
rect 119338 136960 119344 137012
rect 119396 137000 119402 137012
rect 120718 137000 120724 137012
rect 119396 136972 120724 137000
rect 119396 136960 119402 136972
rect 120718 136960 120724 136972
rect 120776 136960 120782 137012
rect 148962 136960 148968 137012
rect 149020 137000 149026 137012
rect 150618 137000 150624 137012
rect 149020 136972 150624 137000
rect 149020 136960 149026 136972
rect 150618 136960 150624 136972
rect 150676 136960 150682 137012
rect 147582 136756 147588 136808
rect 147640 136796 147646 136808
rect 149054 136796 149060 136808
rect 147640 136768 149060 136796
rect 147640 136756 147646 136768
rect 149054 136756 149060 136768
rect 149112 136756 149118 136808
rect 160002 136688 160008 136740
rect 160060 136728 160066 136740
rect 161474 136728 161480 136740
rect 160060 136700 161480 136728
rect 160060 136688 160066 136700
rect 161474 136688 161480 136700
rect 161532 136688 161538 136740
rect 3326 136620 3332 136672
rect 3384 136660 3390 136672
rect 112530 136660 112536 136672
rect 3384 136632 112536 136660
rect 3384 136620 3390 136632
rect 112530 136620 112536 136632
rect 112588 136620 112594 136672
rect 45002 135872 45008 135924
rect 45060 135912 45066 135924
rect 178126 135912 178132 135924
rect 45060 135884 178132 135912
rect 45060 135872 45066 135884
rect 178126 135872 178132 135884
rect 178184 135872 178190 135924
rect 116486 129820 116492 129872
rect 116544 129860 116550 129872
rect 116670 129860 116676 129872
rect 116544 129832 116676 129860
rect 116544 129820 116550 129832
rect 116670 129820 116676 129832
rect 116728 129820 116734 129872
rect 97258 129072 97264 129124
rect 97316 129112 97322 129124
rect 102778 129112 102784 129124
rect 97316 129084 102784 129112
rect 97316 129072 97322 129084
rect 102778 129072 102784 129084
rect 102836 129072 102842 129124
rect 102778 117308 102784 117360
rect 102836 117348 102842 117360
rect 102836 117320 103514 117348
rect 102836 117308 102842 117320
rect 103486 117280 103514 117320
rect 105538 117280 105544 117292
rect 103486 117252 105544 117280
rect 105538 117240 105544 117252
rect 105596 117240 105602 117292
rect 87598 104796 87604 104848
rect 87656 104836 87662 104848
rect 90358 104836 90364 104848
rect 87656 104808 90364 104836
rect 87656 104796 87662 104808
rect 90358 104796 90364 104808
rect 90416 104796 90422 104848
rect 116486 100308 116492 100360
rect 116544 100348 116550 100360
rect 116762 100348 116768 100360
rect 116544 100320 116768 100348
rect 116544 100308 116550 100320
rect 116762 100308 116768 100320
rect 116820 100308 116826 100360
rect 90358 99968 90364 100020
rect 90416 100008 90422 100020
rect 101398 100008 101404 100020
rect 90416 99980 101404 100008
rect 90416 99968 90422 99980
rect 101398 99968 101404 99980
rect 101456 99968 101462 100020
rect 177390 99356 177396 99408
rect 177448 99396 177454 99408
rect 580166 99396 580172 99408
rect 177448 99368 580172 99396
rect 177448 99356 177454 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 105538 92488 105544 92540
rect 105596 92528 105602 92540
rect 109402 92528 109408 92540
rect 105596 92500 109408 92528
rect 105596 92488 105602 92500
rect 109402 92488 109408 92500
rect 109460 92488 109466 92540
rect 109402 89700 109408 89752
rect 109460 89740 109466 89752
rect 109460 89712 113174 89740
rect 109460 89700 109466 89712
rect 101398 89632 101404 89684
rect 101456 89672 101462 89684
rect 104158 89672 104164 89684
rect 101456 89644 104164 89672
rect 101456 89632 101462 89644
rect 104158 89632 104164 89644
rect 104216 89632 104222 89684
rect 113146 89672 113174 89712
rect 114370 89672 114376 89684
rect 113146 89644 114376 89672
rect 114370 89632 114376 89644
rect 114428 89632 114434 89684
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 116670 84232 116676 84244
rect 3384 84204 116676 84232
rect 3384 84192 3390 84204
rect 116670 84192 116676 84204
rect 116728 84192 116734 84244
rect 175274 76508 175280 76560
rect 175332 76548 175338 76560
rect 527174 76548 527180 76560
rect 175332 76520 527180 76548
rect 175332 76508 175338 76520
rect 527174 76508 527180 76520
rect 527232 76508 527238 76560
rect 421558 75868 421564 75880
rect 176626 75840 421564 75868
rect 164206 75772 170536 75800
rect 43622 75692 43628 75744
rect 43680 75732 43686 75744
rect 164206 75732 164234 75772
rect 43680 75704 164234 75732
rect 166966 75704 169754 75732
rect 43680 75692 43686 75704
rect 114554 75624 114560 75676
rect 114612 75664 114618 75676
rect 119982 75664 119988 75676
rect 114612 75636 119988 75664
rect 114612 75624 114618 75636
rect 119982 75624 119988 75636
rect 120040 75624 120046 75676
rect 166966 75664 166994 75704
rect 154040 75636 158714 75664
rect 13078 75556 13084 75608
rect 13136 75596 13142 75608
rect 13136 75568 135484 75596
rect 13136 75556 13142 75568
rect 4890 75488 4896 75540
rect 4948 75528 4954 75540
rect 4948 75500 132494 75528
rect 4948 75488 4954 75500
rect 132466 74712 132494 75500
rect 135456 74792 135484 75568
rect 147646 75364 149054 75392
rect 147646 75256 147674 75364
rect 135640 75228 142154 75256
rect 135438 74740 135444 74792
rect 135496 74740 135502 74792
rect 135640 74712 135668 75228
rect 142126 75188 142154 75228
rect 143506 75228 144914 75256
rect 143506 75188 143534 75228
rect 142126 75160 143534 75188
rect 144886 75188 144914 75228
rect 146266 75228 147674 75256
rect 146266 75188 146294 75228
rect 144886 75160 146294 75188
rect 149026 75188 149054 75364
rect 154040 75188 154068 75636
rect 158686 75596 158714 75636
rect 165586 75636 166994 75664
rect 158686 75568 160094 75596
rect 160066 75528 160094 75568
rect 162826 75568 164234 75596
rect 160066 75500 161474 75528
rect 161446 75460 161474 75500
rect 162826 75460 162854 75568
rect 161446 75432 162854 75460
rect 164206 75460 164234 75568
rect 165586 75460 165614 75636
rect 169726 75528 169754 75704
rect 170508 75676 170536 75772
rect 176626 75732 176654 75840
rect 421558 75828 421564 75840
rect 421616 75828 421622 75880
rect 417418 75800 417424 75812
rect 170600 75704 176654 75732
rect 180766 75772 417424 75800
rect 170600 75676 170628 75704
rect 170490 75624 170496 75676
rect 170548 75624 170554 75676
rect 170582 75624 170588 75676
rect 170640 75624 170646 75676
rect 170674 75624 170680 75676
rect 170732 75664 170738 75676
rect 177390 75664 177396 75676
rect 170732 75636 177396 75664
rect 170732 75624 170738 75636
rect 177390 75624 177396 75636
rect 177448 75624 177454 75676
rect 170398 75528 170404 75540
rect 169726 75500 170404 75528
rect 170398 75488 170404 75500
rect 170456 75488 170462 75540
rect 164206 75432 165614 75460
rect 170674 75284 170680 75336
rect 170732 75324 170738 75336
rect 180766 75324 180794 75772
rect 417418 75760 417424 75772
rect 417476 75760 417482 75812
rect 170732 75296 180794 75324
rect 170732 75284 170738 75296
rect 149026 75160 154068 75188
rect 154132 75228 155908 75256
rect 154132 75120 154160 75228
rect 132466 74684 135668 74712
rect 138400 75092 142154 75120
rect 135438 74536 135444 74588
rect 135496 74576 135502 74588
rect 138400 74576 138428 75092
rect 142126 75052 142154 75092
rect 143506 75092 154160 75120
rect 154546 75092 155724 75120
rect 143506 75052 143534 75092
rect 154546 75052 154574 75092
rect 142126 75024 143534 75052
rect 143644 75024 154574 75052
rect 143644 74780 143672 75024
rect 146312 74956 155356 74984
rect 143718 74876 143724 74928
rect 143776 74916 143782 74928
rect 146312 74916 146340 74956
rect 143776 74888 146340 74916
rect 143776 74876 143782 74888
rect 146478 74876 146484 74928
rect 146536 74876 146542 74928
rect 146496 74848 146524 74876
rect 146496 74820 149836 74848
rect 143718 74780 143724 74792
rect 143644 74752 143724 74780
rect 143718 74740 143724 74752
rect 143776 74740 143782 74792
rect 135496 74548 138428 74576
rect 135496 74536 135502 74548
rect 149808 74508 149836 74820
rect 155328 74576 155356 74956
rect 155696 74644 155724 75092
rect 155880 74712 155908 75228
rect 172422 75216 172428 75268
rect 172480 75256 172486 75268
rect 462314 75256 462320 75268
rect 172480 75228 462320 75256
rect 172480 75216 172486 75228
rect 462314 75216 462320 75228
rect 462372 75216 462378 75268
rect 580258 75188 580264 75200
rect 176626 75160 580264 75188
rect 158548 75092 164234 75120
rect 158548 74984 158576 75092
rect 164206 75052 164234 75092
rect 164206 75024 169754 75052
rect 157720 74956 158576 74984
rect 169726 74984 169754 75024
rect 170674 74984 170680 74996
rect 169726 74956 170680 74984
rect 157720 74792 157748 74956
rect 170674 74944 170680 74956
rect 170732 74944 170738 74996
rect 170950 74944 170956 74996
rect 171008 74984 171014 74996
rect 176626 74984 176654 75160
rect 580258 75148 580264 75160
rect 580316 75148 580322 75200
rect 171008 74956 176654 74984
rect 171008 74944 171014 74956
rect 168374 74876 168380 74928
rect 168432 74916 168438 74928
rect 172422 74916 172428 74928
rect 168432 74888 172428 74916
rect 168432 74876 168438 74888
rect 172422 74876 172428 74888
rect 172480 74876 172486 74928
rect 169570 74848 169576 74860
rect 157812 74820 169576 74848
rect 157702 74740 157708 74792
rect 157760 74740 157766 74792
rect 157812 74712 157840 74820
rect 169570 74808 169576 74820
rect 169628 74808 169634 74860
rect 169754 74808 169760 74860
rect 169812 74848 169818 74860
rect 170490 74848 170496 74860
rect 169812 74820 170496 74848
rect 169812 74808 169818 74820
rect 170490 74808 170496 74820
rect 170548 74808 170554 74860
rect 170674 74808 170680 74860
rect 170732 74848 170738 74860
rect 235810 74848 235816 74860
rect 170732 74820 235816 74848
rect 170732 74808 170738 74820
rect 235810 74808 235816 74820
rect 235868 74808 235874 74860
rect 249978 74780 249984 74792
rect 155880 74684 157840 74712
rect 157904 74752 249984 74780
rect 157904 74644 157932 74752
rect 249978 74740 249984 74752
rect 250036 74740 250042 74792
rect 285398 74712 285404 74724
rect 155696 74616 157932 74644
rect 157996 74684 285404 74712
rect 157996 74576 158024 74684
rect 285398 74672 285404 74684
rect 285456 74672 285462 74724
rect 320910 74644 320916 74656
rect 155328 74548 155448 74576
rect 155420 74508 155448 74548
rect 155604 74548 158024 74576
rect 159652 74616 320916 74644
rect 155604 74508 155632 74548
rect 118666 74480 144914 74508
rect 149808 74480 155356 74508
rect 155420 74480 155632 74508
rect 112530 74332 112536 74384
rect 112588 74372 112594 74384
rect 118666 74372 118694 74480
rect 144886 74372 144914 74480
rect 148226 74400 148232 74452
rect 148284 74440 148290 74452
rect 148284 74412 155172 74440
rect 148284 74400 148290 74412
rect 112588 74344 118694 74372
rect 128326 74344 138014 74372
rect 144886 74344 155080 74372
rect 112588 74332 112594 74344
rect 116670 74264 116676 74316
rect 116728 74304 116734 74316
rect 128326 74304 128354 74344
rect 116728 74276 128354 74304
rect 137986 74304 138014 74344
rect 148226 74304 148232 74316
rect 137986 74276 148232 74304
rect 116728 74264 116734 74276
rect 148226 74264 148232 74276
rect 148284 74264 148290 74316
rect 112438 74196 112444 74248
rect 112496 74236 112502 74248
rect 112496 74208 118694 74236
rect 112496 74196 112502 74208
rect 118666 73896 118694 74208
rect 137986 74208 154988 74236
rect 137986 73896 138014 74208
rect 152274 74128 152280 74180
rect 152332 74168 152338 74180
rect 152734 74168 152740 74180
rect 152332 74140 152740 74168
rect 152332 74128 152338 74140
rect 152734 74128 152740 74140
rect 152792 74128 152798 74180
rect 148226 74060 148232 74112
rect 148284 74100 148290 74112
rect 148284 74072 150434 74100
rect 148284 74060 148290 74072
rect 139578 73924 139584 73976
rect 139636 73964 139642 73976
rect 141418 73964 141424 73976
rect 139636 73936 141424 73964
rect 139636 73924 139642 73936
rect 141418 73924 141424 73936
rect 141476 73924 141482 73976
rect 118666 73868 138014 73896
rect 140774 73788 140780 73840
rect 140832 73828 140838 73840
rect 141418 73828 141424 73840
rect 140832 73800 141424 73828
rect 140832 73788 140838 73800
rect 141418 73788 141424 73800
rect 141476 73788 141482 73840
rect 150406 73828 150434 74072
rect 152734 73924 152740 73976
rect 152792 73964 152798 73976
rect 153102 73964 153108 73976
rect 152792 73936 153108 73964
rect 152792 73924 152798 73936
rect 153102 73924 153108 73936
rect 153160 73924 153166 73976
rect 154960 73964 154988 74208
rect 155052 74032 155080 74344
rect 155144 74100 155172 74412
rect 155328 74372 155356 74480
rect 159652 74440 159680 74616
rect 320910 74604 320916 74616
rect 320968 74604 320974 74656
rect 343358 74576 343364 74588
rect 164206 74548 343364 74576
rect 164206 74440 164234 74548
rect 343358 74536 343364 74548
rect 343416 74536 343422 74588
rect 167730 74468 167736 74520
rect 167788 74508 167794 74520
rect 413278 74508 413284 74520
rect 167788 74480 413284 74508
rect 167788 74468 167794 74480
rect 413278 74468 413284 74480
rect 413336 74468 413342 74520
rect 155512 74412 159680 74440
rect 160066 74412 164234 74440
rect 155512 74372 155540 74412
rect 160066 74372 160094 74412
rect 167454 74400 167460 74452
rect 167512 74440 167518 74452
rect 410518 74440 410524 74452
rect 167512 74412 410524 74440
rect 167512 74400 167518 74412
rect 410518 74400 410524 74412
rect 410576 74400 410582 74452
rect 170030 74372 170036 74384
rect 155328 74344 155540 74372
rect 158824 74344 160094 74372
rect 162826 74344 170036 74372
rect 158824 74168 158852 74344
rect 162826 74304 162854 74344
rect 170030 74332 170036 74344
rect 170088 74332 170094 74384
rect 169938 74304 169944 74316
rect 158732 74140 158852 74168
rect 159008 74276 162854 74304
rect 164206 74276 169944 74304
rect 158732 74100 158760 74140
rect 155144 74072 158760 74100
rect 159008 74032 159036 74276
rect 164206 74236 164234 74276
rect 169938 74264 169944 74276
rect 169996 74264 170002 74316
rect 155052 74004 159036 74032
rect 159100 74208 164234 74236
rect 159100 73964 159128 74208
rect 168466 74196 168472 74248
rect 168524 74236 168530 74248
rect 397454 74236 397460 74248
rect 168524 74208 397460 74236
rect 168524 74196 168530 74208
rect 397454 74196 397460 74208
rect 397512 74196 397518 74248
rect 159174 74128 159180 74180
rect 159232 74168 159238 74180
rect 484026 74168 484032 74180
rect 159232 74140 484032 74168
rect 159232 74128 159238 74140
rect 484026 74128 484032 74140
rect 484084 74128 484090 74180
rect 170122 74100 170128 74112
rect 154960 73936 159128 73964
rect 160066 74072 170128 74100
rect 160066 73828 160094 74072
rect 170122 74060 170128 74072
rect 170180 74060 170186 74112
rect 171778 74060 171784 74112
rect 171836 74100 171842 74112
rect 515950 74100 515956 74112
rect 171836 74072 515956 74100
rect 171836 74060 171842 74072
rect 515950 74060 515956 74072
rect 516008 74060 516014 74112
rect 163038 73992 163044 74044
rect 163096 74032 163102 74044
rect 533706 74032 533712 74044
rect 163096 74004 533712 74032
rect 163096 73992 163102 74004
rect 533706 73992 533712 74004
rect 533764 73992 533770 74044
rect 164418 73924 164424 73976
rect 164476 73964 164482 73976
rect 551462 73964 551468 73976
rect 164476 73936 551468 73964
rect 164476 73924 164482 73936
rect 551462 73924 551468 73936
rect 551520 73924 551526 73976
rect 163314 73856 163320 73908
rect 163372 73896 163378 73908
rect 537202 73896 537208 73908
rect 163372 73868 537208 73896
rect 163372 73856 163378 73868
rect 537202 73856 537208 73868
rect 537260 73856 537266 73908
rect 150406 73800 160094 73828
rect 164694 73788 164700 73840
rect 164752 73828 164758 73840
rect 554958 73828 554964 73840
rect 164752 73800 554964 73828
rect 164752 73788 164758 73800
rect 554958 73788 554964 73800
rect 555016 73788 555022 73840
rect 5074 73720 5080 73772
rect 5132 73760 5138 73772
rect 5132 73732 150434 73760
rect 5132 73720 5138 73732
rect 140958 73652 140964 73704
rect 141016 73692 141022 73704
rect 150406 73692 150434 73732
rect 161658 73720 161664 73772
rect 161716 73760 161722 73772
rect 171778 73760 171784 73772
rect 161716 73732 171784 73760
rect 161716 73720 161722 73732
rect 171778 73720 171784 73732
rect 171836 73720 171842 73772
rect 169662 73692 169668 73704
rect 141016 73664 142108 73692
rect 150406 73664 169668 73692
rect 141016 73652 141022 73664
rect 140774 73584 140780 73636
rect 140832 73624 140838 73636
rect 141050 73624 141056 73636
rect 140832 73596 141056 73624
rect 140832 73584 140838 73596
rect 141050 73584 141056 73596
rect 141108 73584 141114 73636
rect 141694 73584 141700 73636
rect 141752 73584 141758 73636
rect 140958 73448 140964 73500
rect 141016 73488 141022 73500
rect 141234 73488 141240 73500
rect 141016 73460 141240 73488
rect 141016 73448 141022 73460
rect 141234 73448 141240 73460
rect 141292 73448 141298 73500
rect 141142 73380 141148 73432
rect 141200 73420 141206 73432
rect 141510 73420 141516 73432
rect 141200 73392 141516 73420
rect 141200 73380 141206 73392
rect 141510 73380 141516 73392
rect 141568 73380 141574 73432
rect 122926 73312 122932 73364
rect 122984 73352 122990 73364
rect 123662 73352 123668 73364
rect 122984 73324 123668 73352
rect 122984 73312 122990 73324
rect 123662 73312 123668 73324
rect 123720 73312 123726 73364
rect 141234 73312 141240 73364
rect 141292 73352 141298 73364
rect 141712 73352 141740 73584
rect 142080 73432 142108 73664
rect 169662 73652 169668 73664
rect 169720 73652 169726 73704
rect 167914 73584 167920 73636
rect 167972 73624 167978 73636
rect 172698 73624 172704 73636
rect 167972 73596 172704 73624
rect 167972 73584 167978 73596
rect 172698 73584 172704 73596
rect 172756 73584 172762 73636
rect 167638 73516 167644 73568
rect 167696 73556 167702 73568
rect 170582 73556 170588 73568
rect 167696 73528 170588 73556
rect 167696 73516 167702 73528
rect 170582 73516 170588 73528
rect 170640 73516 170646 73568
rect 168098 73448 168104 73500
rect 168156 73488 168162 73500
rect 170950 73488 170956 73500
rect 168156 73460 170956 73488
rect 168156 73448 168162 73460
rect 170950 73448 170956 73460
rect 171008 73448 171014 73500
rect 142062 73380 142068 73432
rect 142120 73380 142126 73432
rect 141292 73324 141740 73352
rect 141292 73312 141298 73324
rect 158898 73312 158904 73364
rect 158956 73352 158962 73364
rect 163038 73352 163044 73364
rect 158956 73324 163044 73352
rect 158956 73312 158962 73324
rect 163038 73312 163044 73324
rect 163096 73312 163102 73364
rect 150360 73256 150572 73284
rect 124306 73216 124312 73228
rect 124140 73188 124312 73216
rect 124140 73148 124168 73188
rect 124306 73176 124312 73188
rect 124364 73176 124370 73228
rect 118666 73120 124168 73148
rect 113910 72768 113916 72820
rect 113968 72808 113974 72820
rect 118666 72808 118694 73120
rect 141418 73108 141424 73160
rect 141476 73148 141482 73160
rect 142338 73148 142344 73160
rect 141476 73120 142344 73148
rect 141476 73108 141482 73120
rect 142338 73108 142344 73120
rect 142396 73108 142402 73160
rect 143074 73108 143080 73160
rect 143132 73148 143138 73160
rect 150360 73148 150388 73256
rect 150434 73176 150440 73228
rect 150492 73176 150498 73228
rect 143132 73120 150388 73148
rect 143132 73108 143138 73120
rect 119614 73040 119620 73092
rect 119672 73080 119678 73092
rect 130378 73080 130384 73092
rect 119672 73052 130384 73080
rect 119672 73040 119678 73052
rect 130378 73040 130384 73052
rect 130436 73040 130442 73092
rect 147766 73040 147772 73092
rect 147824 73080 147830 73092
rect 148226 73080 148232 73092
rect 147824 73052 148232 73080
rect 147824 73040 147830 73052
rect 148226 73040 148232 73052
rect 148284 73040 148290 73092
rect 121178 72972 121184 73024
rect 121236 73012 121242 73024
rect 129274 73012 129280 73024
rect 121236 72984 129280 73012
rect 121236 72972 121242 72984
rect 129274 72972 129280 72984
rect 129332 72972 129338 73024
rect 136634 72972 136640 73024
rect 136692 73012 136698 73024
rect 139854 73012 139860 73024
rect 136692 72984 139860 73012
rect 136692 72972 136698 72984
rect 139854 72972 139860 72984
rect 139912 72972 139918 73024
rect 123110 72904 123116 72956
rect 123168 72944 123174 72956
rect 123570 72944 123576 72956
rect 123168 72916 123576 72944
rect 123168 72904 123174 72916
rect 123570 72904 123576 72916
rect 123628 72904 123634 72956
rect 124324 72916 128354 72944
rect 113968 72780 118694 72808
rect 113968 72768 113974 72780
rect 121270 72768 121276 72820
rect 121328 72808 121334 72820
rect 124324 72808 124352 72916
rect 125226 72836 125232 72888
rect 125284 72836 125290 72888
rect 128326 72876 128354 72916
rect 129734 72904 129740 72956
rect 129792 72944 129798 72956
rect 129918 72944 129924 72956
rect 129792 72916 129924 72944
rect 129792 72904 129798 72916
rect 129918 72904 129924 72916
rect 129976 72904 129982 72956
rect 130378 72904 130384 72956
rect 130436 72944 130442 72956
rect 130562 72944 130568 72956
rect 130436 72916 130568 72944
rect 130436 72904 130442 72916
rect 130562 72904 130568 72916
rect 130620 72904 130626 72956
rect 129826 72876 129832 72888
rect 128326 72848 129832 72876
rect 129826 72836 129832 72848
rect 129884 72836 129890 72888
rect 145098 72836 145104 72888
rect 145156 72876 145162 72888
rect 145156 72848 147674 72876
rect 145156 72836 145162 72848
rect 125244 72808 125272 72836
rect 121328 72780 124352 72808
rect 124600 72780 125272 72808
rect 121328 72768 121334 72780
rect 124600 72752 124628 72780
rect 130286 72768 130292 72820
rect 130344 72808 130350 72820
rect 130562 72808 130568 72820
rect 130344 72780 130568 72808
rect 130344 72768 130350 72780
rect 130562 72768 130568 72780
rect 130620 72768 130626 72820
rect 118142 72700 118148 72752
rect 118200 72740 118206 72752
rect 123754 72740 123760 72752
rect 118200 72712 123760 72740
rect 118200 72700 118206 72712
rect 123754 72700 123760 72712
rect 123812 72700 123818 72752
rect 124582 72700 124588 72752
rect 124640 72700 124646 72752
rect 125226 72700 125232 72752
rect 125284 72740 125290 72752
rect 125502 72740 125508 72752
rect 125284 72712 125508 72740
rect 125284 72700 125290 72712
rect 125502 72700 125508 72712
rect 125560 72700 125566 72752
rect 126422 72700 126428 72752
rect 126480 72740 126486 72752
rect 126790 72740 126796 72752
rect 126480 72712 126796 72740
rect 126480 72700 126486 72712
rect 126790 72700 126796 72712
rect 126848 72700 126854 72752
rect 129918 72700 129924 72752
rect 129976 72740 129982 72752
rect 130102 72740 130108 72752
rect 129976 72712 130108 72740
rect 129976 72700 129982 72712
rect 130102 72700 130108 72712
rect 130160 72700 130166 72752
rect 134610 72700 134616 72752
rect 134668 72740 134674 72752
rect 135070 72740 135076 72752
rect 134668 72712 135076 72740
rect 134668 72700 134674 72712
rect 135070 72700 135076 72712
rect 135128 72700 135134 72752
rect 145098 72700 145104 72752
rect 145156 72740 145162 72752
rect 145834 72740 145840 72752
rect 145156 72712 145840 72740
rect 145156 72700 145162 72712
rect 145834 72700 145840 72712
rect 145892 72700 145898 72752
rect 109678 72632 109684 72684
rect 109736 72672 109742 72684
rect 109736 72644 123156 72672
rect 109736 72632 109742 72644
rect 107010 72496 107016 72548
rect 107068 72536 107074 72548
rect 123018 72536 123024 72548
rect 107068 72508 123024 72536
rect 107068 72496 107074 72508
rect 123018 72496 123024 72508
rect 123076 72496 123082 72548
rect 123128 72536 123156 72644
rect 123386 72632 123392 72684
rect 123444 72632 123450 72684
rect 124858 72672 124864 72684
rect 123496 72644 124864 72672
rect 123202 72564 123208 72616
rect 123260 72604 123266 72616
rect 123404 72604 123432 72632
rect 123260 72576 123432 72604
rect 123260 72564 123266 72576
rect 123496 72536 123524 72644
rect 124858 72632 124864 72644
rect 124916 72632 124922 72684
rect 141602 72632 141608 72684
rect 141660 72672 141666 72684
rect 141786 72672 141792 72684
rect 141660 72644 141792 72672
rect 141660 72632 141666 72644
rect 141786 72632 141792 72644
rect 141844 72632 141850 72684
rect 147646 72672 147674 72848
rect 150452 72808 150480 73176
rect 150544 73148 150572 73256
rect 152274 73244 152280 73296
rect 152332 73284 152338 73296
rect 152332 73256 154574 73284
rect 152332 73244 152338 73256
rect 151354 73176 151360 73228
rect 151412 73216 151418 73228
rect 151412 73188 153792 73216
rect 151412 73176 151418 73188
rect 152274 73148 152280 73160
rect 150544 73120 152280 73148
rect 152274 73108 152280 73120
rect 152332 73108 152338 73160
rect 153286 73108 153292 73160
rect 153344 73148 153350 73160
rect 153344 73120 153516 73148
rect 153344 73108 153350 73120
rect 152366 72972 152372 73024
rect 152424 73012 152430 73024
rect 152424 72984 153148 73012
rect 152424 72972 152430 72984
rect 153120 72888 153148 72984
rect 153102 72836 153108 72888
rect 153160 72836 153166 72888
rect 150452 72780 151676 72808
rect 151648 72752 151676 72780
rect 152366 72768 152372 72820
rect 152424 72808 152430 72820
rect 152642 72808 152648 72820
rect 152424 72780 152648 72808
rect 152424 72768 152430 72780
rect 152642 72768 152648 72780
rect 152700 72768 152706 72820
rect 151078 72700 151084 72752
rect 151136 72740 151142 72752
rect 151354 72740 151360 72752
rect 151136 72712 151360 72740
rect 151136 72700 151142 72712
rect 151354 72700 151360 72712
rect 151412 72700 151418 72752
rect 151630 72700 151636 72752
rect 151688 72700 151694 72752
rect 153488 72740 153516 73120
rect 153764 72944 153792 73188
rect 154546 73012 154574 73256
rect 158806 73244 158812 73296
rect 158864 73284 158870 73296
rect 158864 73256 160784 73284
rect 158864 73244 158870 73256
rect 157978 73176 157984 73228
rect 158036 73176 158042 73228
rect 154942 73108 154948 73160
rect 155000 73148 155006 73160
rect 157702 73148 157708 73160
rect 155000 73120 157708 73148
rect 155000 73108 155006 73120
rect 157702 73108 157708 73120
rect 157760 73108 157766 73160
rect 157996 73148 158024 73176
rect 158806 73148 158812 73160
rect 157996 73120 158812 73148
rect 158806 73108 158812 73120
rect 158864 73108 158870 73160
rect 160756 73148 160784 73256
rect 168374 73244 168380 73296
rect 168432 73284 168438 73296
rect 168834 73284 168840 73296
rect 168432 73256 168840 73284
rect 168432 73244 168438 73256
rect 168834 73244 168840 73256
rect 168892 73244 168898 73296
rect 160830 73176 160836 73228
rect 160888 73216 160894 73228
rect 505370 73216 505376 73228
rect 160888 73188 505376 73216
rect 160888 73176 160894 73188
rect 505370 73176 505376 73188
rect 505428 73176 505434 73228
rect 164418 73148 164424 73160
rect 160756 73120 164424 73148
rect 164418 73108 164424 73120
rect 164476 73108 164482 73160
rect 168282 73108 168288 73160
rect 168340 73148 168346 73160
rect 175274 73148 175280 73160
rect 168340 73120 175280 73148
rect 168340 73108 168346 73120
rect 175274 73108 175280 73120
rect 175332 73108 175338 73160
rect 155494 73040 155500 73092
rect 155552 73080 155558 73092
rect 155552 73052 156000 73080
rect 155552 73040 155558 73052
rect 155972 73012 156000 73052
rect 156046 73040 156052 73092
rect 156104 73080 156110 73092
rect 158898 73080 158904 73092
rect 156104 73052 158904 73080
rect 156104 73040 156110 73052
rect 158898 73040 158904 73052
rect 158956 73040 158962 73092
rect 159174 73040 159180 73092
rect 159232 73080 159238 73092
rect 160002 73080 160008 73092
rect 159232 73052 160008 73080
rect 159232 73040 159238 73052
rect 160002 73040 160008 73052
rect 160060 73040 160066 73092
rect 165706 73040 165712 73092
rect 165764 73080 165770 73092
rect 166902 73080 166908 73092
rect 165764 73052 166908 73080
rect 165764 73040 165770 73052
rect 166902 73040 166908 73052
rect 166960 73040 166966 73092
rect 167822 73040 167828 73092
rect 167880 73080 167886 73092
rect 178678 73080 178684 73092
rect 167880 73052 178684 73080
rect 167880 73040 167886 73052
rect 178678 73040 178684 73052
rect 178736 73040 178742 73092
rect 167546 73012 167552 73024
rect 154546 72984 155724 73012
rect 155972 72984 167552 73012
rect 153764 72916 155632 72944
rect 153838 72768 153844 72820
rect 153896 72808 153902 72820
rect 155494 72808 155500 72820
rect 153896 72780 155500 72808
rect 153896 72768 153902 72780
rect 155494 72768 155500 72780
rect 155552 72768 155558 72820
rect 155604 72808 155632 72916
rect 155696 72876 155724 72984
rect 167546 72972 167552 72984
rect 167604 72972 167610 73024
rect 168006 72972 168012 73024
rect 168064 73012 168070 73024
rect 172146 73012 172152 73024
rect 168064 72984 172152 73012
rect 168064 72972 168070 72984
rect 172146 72972 172152 72984
rect 172204 72972 172210 73024
rect 172330 72972 172336 73024
rect 172388 73012 172394 73024
rect 422938 73012 422944 73024
rect 172388 72984 173894 73012
rect 172388 72972 172394 72984
rect 157150 72904 157156 72956
rect 157208 72944 157214 72956
rect 168926 72944 168932 72956
rect 157208 72916 168932 72944
rect 157208 72904 157214 72916
rect 168926 72904 168932 72916
rect 168984 72904 168990 72956
rect 173866 72944 173894 72984
rect 177408 72984 422944 73012
rect 177408 72944 177436 72984
rect 422938 72972 422944 72984
rect 422996 72972 423002 73024
rect 173866 72916 177436 72944
rect 178678 72904 178684 72956
rect 178736 72944 178742 72956
rect 418798 72944 418804 72956
rect 178736 72916 418804 72944
rect 178736 72904 178742 72916
rect 418798 72904 418804 72916
rect 418856 72904 418862 72956
rect 162578 72876 162584 72888
rect 155696 72848 162584 72876
rect 162578 72836 162584 72848
rect 162636 72836 162642 72888
rect 162688 72848 166994 72876
rect 157518 72808 157524 72820
rect 155604 72780 157524 72808
rect 157518 72768 157524 72780
rect 157576 72768 157582 72820
rect 159450 72768 159456 72820
rect 159508 72808 159514 72820
rect 160002 72808 160008 72820
rect 159508 72780 160008 72808
rect 159508 72768 159514 72780
rect 160002 72768 160008 72780
rect 160060 72768 160066 72820
rect 160278 72768 160284 72820
rect 160336 72808 160342 72820
rect 160738 72808 160744 72820
rect 160336 72780 160744 72808
rect 160336 72768 160342 72780
rect 160738 72768 160744 72780
rect 160796 72768 160802 72820
rect 162688 72808 162716 72848
rect 160848 72780 162716 72808
rect 166966 72808 166994 72848
rect 172698 72836 172704 72888
rect 172756 72876 172762 72888
rect 396718 72876 396724 72888
rect 172756 72848 396724 72876
rect 172756 72836 172762 72848
rect 396718 72836 396724 72848
rect 396776 72836 396782 72888
rect 167730 72808 167736 72820
rect 166966 72780 167736 72808
rect 160848 72740 160876 72780
rect 167730 72768 167736 72780
rect 167788 72768 167794 72820
rect 168466 72768 168472 72820
rect 168524 72808 168530 72820
rect 168742 72808 168748 72820
rect 168524 72780 168748 72808
rect 168524 72768 168530 72780
rect 168742 72768 168748 72780
rect 168800 72768 168806 72820
rect 397546 72808 397552 72820
rect 173866 72780 397552 72808
rect 153488 72712 160876 72740
rect 162578 72700 162584 72752
rect 162636 72740 162642 72752
rect 168098 72740 168104 72752
rect 162636 72712 168104 72740
rect 162636 72700 162642 72712
rect 168098 72700 168104 72712
rect 168156 72700 168162 72752
rect 168558 72700 168564 72752
rect 168616 72740 168622 72752
rect 173866 72740 173894 72780
rect 397546 72768 397552 72780
rect 397604 72768 397610 72820
rect 168616 72712 173894 72740
rect 168616 72700 168622 72712
rect 167638 72672 167644 72684
rect 147646 72644 167644 72672
rect 167638 72632 167644 72644
rect 167696 72632 167702 72684
rect 168190 72632 168196 72684
rect 168248 72672 168254 72684
rect 177298 72672 177304 72684
rect 168248 72644 177304 72672
rect 168248 72632 168254 72644
rect 177298 72632 177304 72644
rect 177356 72632 177362 72684
rect 123570 72564 123576 72616
rect 123628 72604 123634 72616
rect 150434 72604 150440 72616
rect 123628 72576 150440 72604
rect 123628 72564 123634 72576
rect 150434 72564 150440 72576
rect 150492 72564 150498 72616
rect 152642 72564 152648 72616
rect 152700 72604 152706 72616
rect 152918 72604 152924 72616
rect 152700 72576 152924 72604
rect 152700 72564 152706 72576
rect 152918 72564 152924 72576
rect 152976 72564 152982 72616
rect 153102 72564 153108 72616
rect 153160 72604 153166 72616
rect 153160 72576 154620 72604
rect 153160 72564 153166 72576
rect 123128 72508 123524 72536
rect 124306 72496 124312 72548
rect 124364 72536 124370 72548
rect 153838 72536 153844 72548
rect 124364 72508 153844 72536
rect 124364 72496 124370 72508
rect 153838 72496 153844 72508
rect 153896 72496 153902 72548
rect 154592 72536 154620 72576
rect 154666 72564 154672 72616
rect 154724 72604 154730 72616
rect 154850 72604 154856 72616
rect 154724 72576 154856 72604
rect 154724 72564 154730 72576
rect 154850 72564 154856 72576
rect 154908 72564 154914 72616
rect 156138 72564 156144 72616
rect 156196 72604 156202 72616
rect 445018 72604 445024 72616
rect 156196 72576 445024 72604
rect 156196 72564 156202 72576
rect 445018 72564 445024 72576
rect 445076 72564 445082 72616
rect 154592 72508 157288 72536
rect 157260 72480 157288 72508
rect 161842 72496 161848 72548
rect 161900 72536 161906 72548
rect 162578 72536 162584 72548
rect 161900 72508 162584 72536
rect 161900 72496 161906 72508
rect 162578 72496 162584 72508
rect 162636 72496 162642 72548
rect 163406 72496 163412 72548
rect 163464 72536 163470 72548
rect 163590 72536 163596 72548
rect 163464 72508 163596 72536
rect 163464 72496 163470 72508
rect 163590 72496 163596 72508
rect 163648 72496 163654 72548
rect 164418 72496 164424 72548
rect 164476 72536 164482 72548
rect 471238 72536 471244 72548
rect 164476 72508 471244 72536
rect 164476 72496 164482 72508
rect 471238 72496 471244 72508
rect 471296 72496 471302 72548
rect 23014 72428 23020 72480
rect 23072 72468 23078 72480
rect 123294 72468 123300 72480
rect 23072 72440 103514 72468
rect 23072 72428 23078 72440
rect 103486 72400 103514 72440
rect 118666 72440 123300 72468
rect 118666 72400 118694 72440
rect 123294 72428 123300 72440
rect 123352 72428 123358 72480
rect 123386 72428 123392 72480
rect 123444 72468 123450 72480
rect 153286 72468 153292 72480
rect 123444 72440 153292 72468
rect 123444 72428 123450 72440
rect 153286 72428 153292 72440
rect 153344 72428 153350 72480
rect 157242 72428 157248 72480
rect 157300 72428 157306 72480
rect 160830 72428 160836 72480
rect 160888 72468 160894 72480
rect 161382 72468 161388 72480
rect 160888 72440 161388 72468
rect 160888 72428 160894 72440
rect 161382 72428 161388 72440
rect 161440 72428 161446 72480
rect 161934 72428 161940 72480
rect 161992 72468 161998 72480
rect 162670 72468 162676 72480
rect 161992 72440 162676 72468
rect 161992 72428 161998 72440
rect 162670 72428 162676 72440
rect 162728 72428 162734 72480
rect 163130 72428 163136 72480
rect 163188 72468 163194 72480
rect 163958 72468 163964 72480
rect 163188 72440 163964 72468
rect 163188 72428 163194 72440
rect 163958 72428 163964 72440
rect 164016 72428 164022 72480
rect 166810 72428 166816 72480
rect 166868 72468 166874 72480
rect 580258 72468 580264 72480
rect 166868 72440 580264 72468
rect 166868 72428 166874 72440
rect 580258 72428 580264 72440
rect 580316 72428 580322 72480
rect 127894 72400 127900 72412
rect 103486 72372 118694 72400
rect 123312 72372 127900 72400
rect 120994 72292 121000 72344
rect 121052 72332 121058 72344
rect 123312 72332 123340 72372
rect 127894 72360 127900 72372
rect 127952 72360 127958 72412
rect 130102 72360 130108 72412
rect 130160 72400 130166 72412
rect 130654 72400 130660 72412
rect 130160 72372 130660 72400
rect 130160 72360 130166 72372
rect 130654 72360 130660 72372
rect 130712 72360 130718 72412
rect 133046 72360 133052 72412
rect 133104 72400 133110 72412
rect 133598 72400 133604 72412
rect 133104 72372 133604 72400
rect 133104 72360 133110 72372
rect 133598 72360 133604 72372
rect 133656 72360 133662 72412
rect 148226 72360 148232 72412
rect 148284 72400 148290 72412
rect 148594 72400 148600 72412
rect 148284 72372 148600 72400
rect 148284 72360 148290 72372
rect 148594 72360 148600 72372
rect 148652 72360 148658 72412
rect 152182 72360 152188 72412
rect 152240 72400 152246 72412
rect 152240 72372 154804 72400
rect 152240 72360 152246 72372
rect 121052 72304 123340 72332
rect 121052 72292 121058 72304
rect 123386 72292 123392 72344
rect 123444 72332 123450 72344
rect 124122 72332 124128 72344
rect 123444 72304 124128 72332
rect 123444 72292 123450 72304
rect 124122 72292 124128 72304
rect 124180 72292 124186 72344
rect 128170 72332 128176 72344
rect 124232 72304 128176 72332
rect 120902 72224 120908 72276
rect 120960 72264 120966 72276
rect 124232 72264 124260 72304
rect 128170 72292 128176 72304
rect 128228 72292 128234 72344
rect 132586 72292 132592 72344
rect 132644 72332 132650 72344
rect 133506 72332 133512 72344
rect 132644 72304 133512 72332
rect 132644 72292 132650 72304
rect 133506 72292 133512 72304
rect 133564 72292 133570 72344
rect 135898 72292 135904 72344
rect 135956 72332 135962 72344
rect 136266 72332 136272 72344
rect 135956 72304 136272 72332
rect 135956 72292 135962 72304
rect 136266 72292 136272 72304
rect 136324 72292 136330 72344
rect 149698 72292 149704 72344
rect 149756 72332 149762 72344
rect 153286 72332 153292 72344
rect 149756 72304 153292 72332
rect 149756 72292 149762 72304
rect 153286 72292 153292 72304
rect 153344 72292 153350 72344
rect 120960 72236 124260 72264
rect 120960 72224 120966 72236
rect 124398 72224 124404 72276
rect 124456 72264 124462 72276
rect 126238 72264 126244 72276
rect 124456 72236 126244 72264
rect 124456 72224 124462 72236
rect 126238 72224 126244 72236
rect 126296 72224 126302 72276
rect 150250 72224 150256 72276
rect 150308 72264 150314 72276
rect 152182 72264 152188 72276
rect 150308 72236 152188 72264
rect 150308 72224 150314 72236
rect 152182 72224 152188 72236
rect 152240 72224 152246 72276
rect 124122 72156 124128 72208
rect 124180 72196 124186 72208
rect 126698 72196 126704 72208
rect 124180 72168 126704 72196
rect 124180 72156 124186 72168
rect 126698 72156 126704 72168
rect 126756 72156 126762 72208
rect 127434 72156 127440 72208
rect 127492 72196 127498 72208
rect 127802 72196 127808 72208
rect 127492 72168 127808 72196
rect 127492 72156 127498 72168
rect 127802 72156 127808 72168
rect 127860 72156 127866 72208
rect 149146 72156 149152 72208
rect 149204 72196 149210 72208
rect 154482 72196 154488 72208
rect 149204 72168 154488 72196
rect 149204 72156 149210 72168
rect 154482 72156 154488 72168
rect 154540 72156 154546 72208
rect 123570 72088 123576 72140
rect 123628 72128 123634 72140
rect 125962 72128 125968 72140
rect 123628 72100 125968 72128
rect 123628 72088 123634 72100
rect 125962 72088 125968 72100
rect 126020 72088 126026 72140
rect 135438 72088 135444 72140
rect 135496 72128 135502 72140
rect 135622 72128 135628 72140
rect 135496 72100 135628 72128
rect 135496 72088 135502 72100
rect 135622 72088 135628 72100
rect 135680 72088 135686 72140
rect 138106 72088 138112 72140
rect 138164 72128 138170 72140
rect 139302 72128 139308 72140
rect 138164 72100 139308 72128
rect 138164 72088 138170 72100
rect 139302 72088 139308 72100
rect 139360 72088 139366 72140
rect 154776 72128 154804 72372
rect 157702 72360 157708 72412
rect 157760 72400 157766 72412
rect 168190 72400 168196 72412
rect 157760 72372 168196 72400
rect 157760 72360 157766 72372
rect 168190 72360 168196 72372
rect 168248 72360 168254 72412
rect 156598 72292 156604 72344
rect 156656 72332 156662 72344
rect 169110 72332 169116 72344
rect 156656 72304 169116 72332
rect 156656 72292 156662 72304
rect 169110 72292 169116 72304
rect 169168 72292 169174 72344
rect 156138 72224 156144 72276
rect 156196 72264 156202 72276
rect 158622 72264 158628 72276
rect 156196 72236 158628 72264
rect 156196 72224 156202 72236
rect 158622 72224 158628 72236
rect 158680 72224 158686 72276
rect 160922 72224 160928 72276
rect 160980 72264 160986 72276
rect 161198 72264 161204 72276
rect 160980 72236 161204 72264
rect 160980 72224 160986 72236
rect 161198 72224 161204 72236
rect 161256 72224 161262 72276
rect 155494 72156 155500 72208
rect 155552 72196 155558 72208
rect 161934 72196 161940 72208
rect 155552 72168 161940 72196
rect 155552 72156 155558 72168
rect 161934 72156 161940 72168
rect 161992 72156 161998 72208
rect 163038 72156 163044 72208
rect 163096 72196 163102 72208
rect 169202 72196 169208 72208
rect 163096 72168 169208 72196
rect 163096 72156 163102 72168
rect 169202 72156 169208 72168
rect 169260 72156 169266 72208
rect 158254 72128 158260 72140
rect 154776 72100 158260 72128
rect 158254 72088 158260 72100
rect 158312 72088 158318 72140
rect 167362 72088 167368 72140
rect 167420 72128 167426 72140
rect 580810 72128 580816 72140
rect 167420 72100 580816 72128
rect 167420 72088 167426 72100
rect 580810 72088 580816 72100
rect 580868 72088 580874 72140
rect 119338 72020 119344 72072
rect 119396 72060 119402 72072
rect 129734 72060 129740 72072
rect 119396 72032 129740 72060
rect 119396 72020 119402 72032
rect 129734 72020 129740 72032
rect 129792 72020 129798 72072
rect 132678 72020 132684 72072
rect 132736 72060 132742 72072
rect 134518 72060 134524 72072
rect 132736 72032 134524 72060
rect 132736 72020 132742 72032
rect 134518 72020 134524 72032
rect 134576 72020 134582 72072
rect 160370 72020 160376 72072
rect 160428 72060 160434 72072
rect 160922 72060 160928 72072
rect 160428 72032 160928 72060
rect 160428 72020 160434 72032
rect 160922 72020 160928 72032
rect 160980 72020 160986 72072
rect 164602 72020 164608 72072
rect 164660 72060 164666 72072
rect 165154 72060 165160 72072
rect 164660 72032 165160 72060
rect 164660 72020 164666 72032
rect 165154 72020 165160 72032
rect 165212 72020 165218 72072
rect 166994 72020 167000 72072
rect 167052 72060 167058 72072
rect 580166 72060 580172 72072
rect 167052 72032 580172 72060
rect 167052 72020 167058 72032
rect 580166 72020 580172 72032
rect 580224 72020 580230 72072
rect 122834 71952 122840 72004
rect 122892 71992 122898 72004
rect 131114 71992 131120 72004
rect 122892 71964 131120 71992
rect 122892 71952 122898 71964
rect 131114 71952 131120 71964
rect 131172 71952 131178 72004
rect 154390 71952 154396 72004
rect 154448 71992 154454 72004
rect 167914 71992 167920 72004
rect 154448 71964 167920 71992
rect 154448 71952 154454 71964
rect 167914 71952 167920 71964
rect 167972 71952 167978 72004
rect 120718 71884 120724 71936
rect 120776 71924 120782 71936
rect 126974 71924 126980 71936
rect 120776 71896 126980 71924
rect 120776 71884 120782 71896
rect 126974 71884 126980 71896
rect 127032 71884 127038 71936
rect 151906 71884 151912 71936
rect 151964 71924 151970 71936
rect 151964 71896 157104 71924
rect 151964 71884 151970 71896
rect 116762 71816 116768 71868
rect 116820 71856 116826 71868
rect 123202 71856 123208 71868
rect 116820 71828 123208 71856
rect 116820 71816 116826 71828
rect 123202 71816 123208 71828
rect 123260 71816 123266 71868
rect 127710 71816 127716 71868
rect 127768 71856 127774 71868
rect 131022 71856 131028 71868
rect 127768 71828 131028 71856
rect 127768 71816 127774 71828
rect 131022 71816 131028 71828
rect 131080 71816 131086 71868
rect 149054 71816 149060 71868
rect 149112 71856 149118 71868
rect 149112 71828 155448 71856
rect 149112 71816 149118 71828
rect 118050 71748 118056 71800
rect 118108 71788 118114 71800
rect 122926 71788 122932 71800
rect 118108 71760 122932 71788
rect 118108 71748 118114 71760
rect 122926 71748 122932 71760
rect 122984 71748 122990 71800
rect 128170 71748 128176 71800
rect 128228 71788 128234 71800
rect 131482 71788 131488 71800
rect 128228 71760 131488 71788
rect 128228 71748 128234 71760
rect 131482 71748 131488 71760
rect 131540 71748 131546 71800
rect 146018 71748 146024 71800
rect 146076 71788 146082 71800
rect 149698 71788 149704 71800
rect 146076 71760 149704 71788
rect 146076 71748 146082 71760
rect 149698 71748 149704 71760
rect 149756 71748 149762 71800
rect 155420 71788 155448 71828
rect 155420 71760 155540 71788
rect 155512 71732 155540 71760
rect 156322 71748 156328 71800
rect 156380 71788 156386 71800
rect 156874 71788 156880 71800
rect 156380 71760 156880 71788
rect 156380 71748 156386 71760
rect 156874 71748 156880 71760
rect 156932 71748 156938 71800
rect 157076 71788 157104 71896
rect 158898 71884 158904 71936
rect 158956 71924 158962 71936
rect 168006 71924 168012 71936
rect 158956 71896 168012 71924
rect 158956 71884 158962 71896
rect 168006 71884 168012 71896
rect 168064 71884 168070 71936
rect 157518 71816 157524 71868
rect 157576 71856 157582 71868
rect 157576 71828 158944 71856
rect 157576 71816 157582 71828
rect 158916 71800 158944 71828
rect 161934 71816 161940 71868
rect 161992 71856 161998 71868
rect 167822 71856 167828 71868
rect 161992 71828 167828 71856
rect 161992 71816 161998 71828
rect 167822 71816 167828 71828
rect 167880 71816 167886 71868
rect 157702 71788 157708 71800
rect 157076 71760 157708 71788
rect 157702 71748 157708 71760
rect 157760 71748 157766 71800
rect 158898 71748 158904 71800
rect 158956 71748 158962 71800
rect 160738 71748 160744 71800
rect 160796 71788 160802 71800
rect 165614 71788 165620 71800
rect 160796 71760 165620 71788
rect 160796 71748 160802 71760
rect 165614 71748 165620 71760
rect 165672 71748 165678 71800
rect 119430 71680 119436 71732
rect 119488 71720 119494 71732
rect 122742 71720 122748 71732
rect 119488 71692 122748 71720
rect 119488 71680 119494 71692
rect 122742 71680 122748 71692
rect 122800 71680 122806 71732
rect 155494 71680 155500 71732
rect 155552 71680 155558 71732
rect 165706 71680 165712 71732
rect 165764 71720 165770 71732
rect 171778 71720 171784 71732
rect 165764 71692 171784 71720
rect 165764 71680 165770 71692
rect 171778 71680 171784 71692
rect 171836 71680 171842 71732
rect 171870 71680 171876 71732
rect 171928 71720 171934 71732
rect 580442 71720 580448 71732
rect 171928 71692 580448 71720
rect 171928 71680 171934 71692
rect 580442 71680 580448 71692
rect 580500 71680 580506 71732
rect 120810 71612 120816 71664
rect 120868 71652 120874 71664
rect 126422 71652 126428 71664
rect 120868 71624 126428 71652
rect 120868 71612 120874 71624
rect 126422 71612 126428 71624
rect 126480 71612 126486 71664
rect 140774 71612 140780 71664
rect 140832 71652 140838 71664
rect 251174 71652 251180 71664
rect 140832 71624 251180 71652
rect 140832 71612 140838 71624
rect 251174 71612 251180 71624
rect 251232 71612 251238 71664
rect 117958 71544 117964 71596
rect 118016 71584 118022 71596
rect 124766 71584 124772 71596
rect 118016 71556 124772 71584
rect 118016 71544 118022 71556
rect 124766 71544 124772 71556
rect 124824 71544 124830 71596
rect 140958 71544 140964 71596
rect 141016 71584 141022 71596
rect 253474 71584 253480 71596
rect 141016 71556 253480 71584
rect 141016 71544 141022 71556
rect 253474 71544 253480 71556
rect 253532 71544 253538 71596
rect 143534 71476 143540 71528
rect 143592 71516 143598 71528
rect 283098 71516 283104 71528
rect 143592 71488 283104 71516
rect 143592 71476 143598 71488
rect 283098 71476 283104 71488
rect 283156 71476 283162 71528
rect 143994 71408 144000 71460
rect 144052 71448 144058 71460
rect 288986 71448 288992 71460
rect 144052 71420 288992 71448
rect 144052 71408 144058 71420
rect 288986 71408 288992 71420
rect 289044 71408 289050 71460
rect 145466 71340 145472 71392
rect 145524 71380 145530 71392
rect 307938 71380 307944 71392
rect 145524 71352 307944 71380
rect 145524 71340 145530 71352
rect 307938 71340 307944 71352
rect 307996 71340 308002 71392
rect 121086 71272 121092 71324
rect 121144 71312 121150 71324
rect 130930 71312 130936 71324
rect 121144 71284 130936 71312
rect 121144 71272 121150 71284
rect 130930 71272 130936 71284
rect 130988 71272 130994 71324
rect 151998 71272 152004 71324
rect 152056 71312 152062 71324
rect 391842 71312 391848 71324
rect 152056 71284 391848 71312
rect 152056 71272 152062 71284
rect 391842 71272 391848 71284
rect 391900 71272 391906 71324
rect 111058 71204 111064 71256
rect 111116 71244 111122 71256
rect 129182 71244 129188 71256
rect 111116 71216 129188 71244
rect 111116 71204 111122 71216
rect 129182 71204 129188 71216
rect 129240 71204 129246 71256
rect 448606 71244 448612 71256
rect 157306 71216 448612 71244
rect 84470 71136 84476 71188
rect 84528 71176 84534 71188
rect 128078 71176 128084 71188
rect 84528 71148 128084 71176
rect 84528 71136 84534 71148
rect 128078 71136 128084 71148
rect 128136 71136 128142 71188
rect 156414 71136 156420 71188
rect 156472 71176 156478 71188
rect 157306 71176 157334 71216
rect 448606 71204 448612 71216
rect 448664 71204 448670 71256
rect 156472 71148 157334 71176
rect 156472 71136 156478 71148
rect 161382 71136 161388 71188
rect 161440 71176 161446 71188
rect 504174 71176 504180 71188
rect 161440 71148 504180 71176
rect 161440 71136 161446 71148
rect 504174 71136 504180 71148
rect 504232 71136 504238 71188
rect 41874 71068 41880 71120
rect 41932 71108 41938 71120
rect 117958 71108 117964 71120
rect 41932 71080 117964 71108
rect 41932 71068 41938 71080
rect 117958 71068 117964 71080
rect 118016 71068 118022 71120
rect 167730 71068 167736 71120
rect 167788 71108 167794 71120
rect 168190 71108 168196 71120
rect 167788 71080 168196 71108
rect 167788 71068 167794 71080
rect 168190 71068 168196 71080
rect 168248 71068 168254 71120
rect 171778 71068 171784 71120
rect 171836 71108 171842 71120
rect 538398 71108 538404 71120
rect 171836 71080 538404 71108
rect 171836 71068 171842 71080
rect 538398 71068 538404 71080
rect 538456 71068 538462 71120
rect 29638 71000 29644 71052
rect 29696 71040 29702 71052
rect 29696 71012 103514 71040
rect 29696 71000 29702 71012
rect 103486 70904 103514 71012
rect 142338 71000 142344 71052
rect 142396 71040 142402 71052
rect 142396 71012 147674 71040
rect 142396 71000 142402 71012
rect 139854 70932 139860 70984
rect 139912 70972 139918 70984
rect 147646 70972 147674 71012
rect 164142 71000 164148 71052
rect 164200 71040 164206 71052
rect 545482 71040 545488 71052
rect 164200 71012 545488 71040
rect 164200 71000 164206 71012
rect 545482 71000 545488 71012
rect 545540 71000 545546 71052
rect 247586 70972 247592 70984
rect 139912 70944 145972 70972
rect 147646 70944 247592 70972
rect 139912 70932 139918 70944
rect 123754 70904 123760 70916
rect 103486 70876 123760 70904
rect 123754 70864 123760 70876
rect 123812 70864 123818 70916
rect 145558 70864 145564 70916
rect 145616 70904 145622 70916
rect 145834 70904 145840 70916
rect 145616 70876 145840 70904
rect 145616 70864 145622 70876
rect 145834 70864 145840 70876
rect 145892 70864 145898 70916
rect 145944 70904 145972 70944
rect 247586 70932 247592 70944
rect 247644 70932 247650 70984
rect 194410 70904 194416 70916
rect 145944 70876 194416 70904
rect 194410 70864 194416 70876
rect 194468 70864 194474 70916
rect 136082 70796 136088 70848
rect 136140 70836 136146 70848
rect 170398 70836 170404 70848
rect 136140 70808 170404 70836
rect 136140 70796 136146 70808
rect 170398 70796 170404 70808
rect 170456 70796 170462 70848
rect 116394 70728 116400 70780
rect 116452 70768 116458 70780
rect 130378 70768 130384 70780
rect 116452 70740 130384 70768
rect 116452 70728 116458 70740
rect 130378 70728 130384 70740
rect 130436 70728 130442 70780
rect 167086 70728 167092 70780
rect 167144 70768 167150 70780
rect 171870 70768 171876 70780
rect 167144 70740 171876 70768
rect 167144 70728 167150 70740
rect 171870 70728 171876 70740
rect 171928 70728 171934 70780
rect 157978 70660 157984 70712
rect 158036 70700 158042 70712
rect 167730 70700 167736 70712
rect 158036 70672 167736 70700
rect 158036 70660 158042 70672
rect 167730 70660 167736 70672
rect 167788 70660 167794 70712
rect 130378 70456 130384 70508
rect 130436 70496 130442 70508
rect 131206 70496 131212 70508
rect 130436 70468 131212 70496
rect 130436 70456 130442 70468
rect 131206 70456 131212 70468
rect 131264 70456 131270 70508
rect 121730 70388 121736 70440
rect 121788 70428 121794 70440
rect 122098 70428 122104 70440
rect 121788 70400 122104 70428
rect 121788 70388 121794 70400
rect 122098 70388 122104 70400
rect 122156 70388 122162 70440
rect 161492 70400 162808 70428
rect 3510 70320 3516 70372
rect 3568 70360 3574 70372
rect 161492 70360 161520 70400
rect 3568 70332 161520 70360
rect 162780 70360 162808 70400
rect 169386 70360 169392 70372
rect 162780 70332 169392 70360
rect 3568 70320 3574 70332
rect 169386 70320 169392 70332
rect 169444 70320 169450 70372
rect 43530 70252 43536 70304
rect 43588 70292 43594 70304
rect 162210 70292 162216 70304
rect 43588 70264 162216 70292
rect 43588 70252 43594 70264
rect 162210 70252 162216 70264
rect 162268 70252 162274 70304
rect 145742 70184 145748 70236
rect 145800 70224 145806 70236
rect 311434 70224 311440 70236
rect 145800 70196 311440 70224
rect 145800 70184 145806 70196
rect 311434 70184 311440 70196
rect 311492 70184 311498 70236
rect 134702 70116 134708 70168
rect 134760 70156 134766 70168
rect 134760 70128 138014 70156
rect 134760 70116 134766 70128
rect 118786 69980 118792 70032
rect 118844 70020 118850 70032
rect 130746 70020 130752 70032
rect 118844 69992 130752 70020
rect 118844 69980 118850 69992
rect 130746 69980 130752 69992
rect 130804 69980 130810 70032
rect 80882 69844 80888 69896
rect 80940 69884 80946 69896
rect 127434 69884 127440 69896
rect 80940 69856 127440 69884
rect 80940 69844 80946 69856
rect 127434 69844 127440 69856
rect 127492 69844 127498 69896
rect 71038 69776 71044 69828
rect 71096 69816 71102 69828
rect 126882 69816 126888 69828
rect 71096 69788 126888 69816
rect 71096 69776 71102 69788
rect 126882 69776 126888 69788
rect 126940 69776 126946 69828
rect 54938 69708 54944 69760
rect 54996 69748 55002 69760
rect 125778 69748 125784 69760
rect 54996 69720 125784 69748
rect 54996 69708 55002 69720
rect 125778 69708 125784 69720
rect 125836 69708 125842 69760
rect 47854 69640 47860 69692
rect 47912 69680 47918 69692
rect 124214 69680 124220 69692
rect 47912 69652 124220 69680
rect 47912 69640 47918 69652
rect 124214 69640 124220 69652
rect 124272 69640 124278 69692
rect 137986 69544 138014 70128
rect 155494 70116 155500 70168
rect 155552 70156 155558 70168
rect 354030 70156 354036 70168
rect 155552 70128 354036 70156
rect 155552 70116 155558 70128
rect 354030 70116 354036 70128
rect 354088 70116 354094 70168
rect 151262 70048 151268 70100
rect 151320 70088 151326 70100
rect 382366 70088 382372 70100
rect 151320 70060 382372 70088
rect 151320 70048 151326 70060
rect 382366 70048 382372 70060
rect 382424 70048 382430 70100
rect 157242 69980 157248 70032
rect 157300 70020 157306 70032
rect 396534 70020 396540 70032
rect 157300 69992 396540 70020
rect 157300 69980 157306 69992
rect 396534 69980 396540 69992
rect 396592 69980 396598 70032
rect 153194 69912 153200 69964
rect 153252 69952 153258 69964
rect 153252 69924 157334 69952
rect 153252 69912 153258 69924
rect 157306 69884 157334 69924
rect 161934 69912 161940 69964
rect 161992 69952 161998 69964
rect 403618 69952 403624 69964
rect 161992 69924 403624 69952
rect 161992 69912 161998 69924
rect 403618 69912 403624 69924
rect 403676 69912 403682 69964
rect 407206 69884 407212 69896
rect 157306 69856 407212 69884
rect 407206 69844 407212 69856
rect 407264 69844 407270 69896
rect 157794 69776 157800 69828
rect 157852 69816 157858 69828
rect 466270 69816 466276 69828
rect 157852 69788 466276 69816
rect 157852 69776 157858 69788
rect 466270 69776 466276 69788
rect 466328 69776 466334 69828
rect 158070 69708 158076 69760
rect 158128 69748 158134 69760
rect 469858 69748 469864 69760
rect 158128 69720 469864 69748
rect 158128 69708 158134 69720
rect 469858 69708 469864 69720
rect 469916 69708 469922 69760
rect 160186 69640 160192 69692
rect 160244 69680 160250 69692
rect 497090 69680 497096 69692
rect 160244 69652 497096 69680
rect 160244 69640 160250 69652
rect 497090 69640 497096 69652
rect 497148 69640 497154 69692
rect 148502 69572 148508 69624
rect 148560 69612 148566 69624
rect 189810 69612 189816 69624
rect 148560 69584 189816 69612
rect 148560 69572 148566 69584
rect 189810 69572 189816 69584
rect 189868 69572 189874 69624
rect 137986 69516 166994 69544
rect 116578 69436 116584 69488
rect 116636 69476 116642 69488
rect 116636 69448 162164 69476
rect 116636 69436 116642 69448
rect 152642 69164 152648 69216
rect 152700 69204 152706 69216
rect 161934 69204 161940 69216
rect 152700 69176 161940 69204
rect 152700 69164 152706 69176
rect 161934 69164 161940 69176
rect 161992 69164 161998 69216
rect 162136 69204 162164 69448
rect 166966 69340 166994 69516
rect 169570 69340 169576 69352
rect 166966 69312 169576 69340
rect 169570 69300 169576 69312
rect 169628 69300 169634 69352
rect 162210 69232 162216 69284
rect 162268 69272 162274 69284
rect 169294 69272 169300 69284
rect 162268 69244 169300 69272
rect 162268 69232 162274 69244
rect 169294 69232 169300 69244
rect 169352 69232 169358 69284
rect 168466 69204 168472 69216
rect 162136 69176 168472 69204
rect 168466 69164 168472 69176
rect 168524 69164 168530 69216
rect 119522 69028 119528 69080
rect 119580 69068 119586 69080
rect 125226 69068 125232 69080
rect 119580 69040 125232 69068
rect 119580 69028 119586 69040
rect 125226 69028 125232 69040
rect 125284 69028 125290 69080
rect 134610 68824 134616 68876
rect 134668 68864 134674 68876
rect 167178 68864 167184 68876
rect 134668 68836 167184 68864
rect 134668 68824 134674 68836
rect 167178 68824 167184 68836
rect 167236 68824 167242 68876
rect 135438 68756 135444 68808
rect 135496 68796 135502 68808
rect 181438 68796 181444 68808
rect 135496 68768 181444 68796
rect 135496 68756 135502 68768
rect 181438 68756 181444 68768
rect 181496 68756 181502 68808
rect 117590 68688 117596 68740
rect 117648 68728 117654 68740
rect 130102 68728 130108 68740
rect 117648 68700 130108 68728
rect 117648 68688 117654 68700
rect 130102 68688 130108 68700
rect 130160 68688 130166 68740
rect 139302 68688 139308 68740
rect 139360 68728 139366 68740
rect 213362 68728 213368 68740
rect 139360 68700 213368 68728
rect 139360 68688 139366 68700
rect 213362 68688 213368 68700
rect 213420 68688 213426 68740
rect 113818 68620 113824 68672
rect 113876 68660 113882 68672
rect 130194 68660 130200 68672
rect 113876 68632 130200 68660
rect 113876 68620 113882 68632
rect 130194 68620 130200 68632
rect 130252 68620 130258 68672
rect 140314 68620 140320 68672
rect 140372 68660 140378 68672
rect 241698 68660 241704 68672
rect 140372 68632 241704 68660
rect 140372 68620 140378 68632
rect 241698 68620 241704 68632
rect 241756 68620 241762 68672
rect 105538 68552 105544 68604
rect 105596 68592 105602 68604
rect 129642 68592 129648 68604
rect 105596 68564 129648 68592
rect 105596 68552 105602 68564
rect 129642 68552 129648 68564
rect 129700 68552 129706 68604
rect 157426 68552 157432 68604
rect 157484 68592 157490 68604
rect 461578 68592 461584 68604
rect 157484 68564 461584 68592
rect 157484 68552 157490 68564
rect 461578 68552 461584 68564
rect 461636 68552 461642 68604
rect 93946 68484 93952 68536
rect 94004 68524 94010 68536
rect 128814 68524 128820 68536
rect 94004 68496 128820 68524
rect 94004 68484 94010 68496
rect 128814 68484 128820 68496
rect 128872 68484 128878 68536
rect 164694 68484 164700 68536
rect 164752 68524 164758 68536
rect 553762 68524 553768 68536
rect 164752 68496 553768 68524
rect 164752 68484 164758 68496
rect 553762 68484 553768 68496
rect 553820 68484 553826 68536
rect 58434 68416 58440 68468
rect 58492 68456 58498 68468
rect 126054 68456 126060 68468
rect 58492 68428 126060 68456
rect 58492 68416 58498 68428
rect 126054 68416 126060 68428
rect 126112 68416 126118 68468
rect 133138 68416 133144 68468
rect 133196 68456 133202 68468
rect 135898 68456 135904 68468
rect 133196 68428 135904 68456
rect 133196 68416 133202 68428
rect 135898 68416 135904 68428
rect 135956 68416 135962 68468
rect 164602 68416 164608 68468
rect 164660 68456 164666 68468
rect 560846 68456 560852 68468
rect 164660 68428 560852 68456
rect 164660 68416 164666 68428
rect 560846 68416 560852 68428
rect 560904 68416 560910 68468
rect 30098 68348 30104 68400
rect 30156 68388 30162 68400
rect 123846 68388 123852 68400
rect 30156 68360 123852 68388
rect 30156 68348 30162 68360
rect 123846 68348 123852 68360
rect 123904 68348 123910 68400
rect 166902 68348 166908 68400
rect 166960 68388 166966 68400
rect 568022 68388 568028 68400
rect 166960 68360 568028 68388
rect 166960 68348 166966 68360
rect 568022 68348 568028 68360
rect 568080 68348 568086 68400
rect 7650 68280 7656 68332
rect 7708 68320 7714 68332
rect 121730 68320 121736 68332
rect 7708 68292 121736 68320
rect 7708 68280 7714 68292
rect 121730 68280 121736 68292
rect 121788 68280 121794 68332
rect 166258 68280 166264 68332
rect 166316 68320 166322 68332
rect 575106 68320 575112 68332
rect 166316 68292 575112 68320
rect 166316 68280 166322 68292
rect 575106 68280 575112 68292
rect 575164 68280 575170 68332
rect 141050 68076 141056 68128
rect 141108 68116 141114 68128
rect 141510 68116 141516 68128
rect 141108 68088 141516 68116
rect 141108 68076 141114 68088
rect 141510 68076 141516 68088
rect 141568 68076 141574 68128
rect 130470 67600 130476 67652
rect 130528 67640 130534 67652
rect 131390 67640 131396 67652
rect 130528 67612 131396 67640
rect 130528 67600 130534 67612
rect 131390 67600 131396 67612
rect 131448 67600 131454 67652
rect 150802 67532 150808 67584
rect 150860 67572 150866 67584
rect 151538 67572 151544 67584
rect 150860 67544 151544 67572
rect 150860 67532 150866 67544
rect 151538 67532 151544 67544
rect 151596 67532 151602 67584
rect 142798 67464 142804 67516
rect 142856 67504 142862 67516
rect 143074 67504 143080 67516
rect 142856 67476 143080 67504
rect 142856 67464 142862 67476
rect 143074 67464 143080 67476
rect 143132 67464 143138 67516
rect 155954 67464 155960 67516
rect 156012 67504 156018 67516
rect 156782 67504 156788 67516
rect 156012 67476 156788 67504
rect 156012 67464 156018 67476
rect 156782 67464 156788 67476
rect 156840 67464 156846 67516
rect 115198 67124 115204 67176
rect 115256 67164 115262 67176
rect 130286 67164 130292 67176
rect 115256 67136 130292 67164
rect 115256 67124 115262 67136
rect 130286 67124 130292 67136
rect 130344 67124 130350 67176
rect 161290 67124 161296 67176
rect 161348 67164 161354 67176
rect 170582 67164 170588 67176
rect 161348 67136 170588 67164
rect 161348 67124 161354 67136
rect 170582 67124 170588 67136
rect 170640 67124 170646 67176
rect 103330 67056 103336 67108
rect 103388 67096 103394 67108
rect 129550 67096 129556 67108
rect 103388 67068 129556 67096
rect 103388 67056 103394 67068
rect 129550 67056 129556 67068
rect 129608 67056 129614 67108
rect 146938 67056 146944 67108
rect 146996 67096 147002 67108
rect 326798 67096 326804 67108
rect 146996 67068 326804 67096
rect 146996 67056 147002 67068
rect 326798 67056 326804 67068
rect 326856 67056 326862 67108
rect 332594 67056 332600 67108
rect 332652 67096 332658 67108
rect 472250 67096 472256 67108
rect 332652 67068 472256 67096
rect 332652 67056 332658 67068
rect 472250 67056 472256 67068
rect 472308 67056 472314 67108
rect 97442 66988 97448 67040
rect 97500 67028 97506 67040
rect 129090 67028 129096 67040
rect 97500 67000 129096 67028
rect 97500 66988 97506 67000
rect 129090 66988 129096 67000
rect 129148 66988 129154 67040
rect 141234 66988 141240 67040
rect 141292 67028 141298 67040
rect 141694 67028 141700 67040
rect 141292 67000 141700 67028
rect 141292 66988 141298 67000
rect 141694 66988 141700 67000
rect 141752 66988 141758 67040
rect 148870 66988 148876 67040
rect 148928 67028 148934 67040
rect 348050 67028 348056 67040
rect 148928 67000 348056 67028
rect 148928 66988 148934 67000
rect 348050 66988 348056 67000
rect 348108 66988 348114 67040
rect 76190 66920 76196 66972
rect 76248 66960 76254 66972
rect 127066 66960 127072 66972
rect 76248 66932 127072 66960
rect 76248 66920 76254 66932
rect 127066 66920 127072 66932
rect 127124 66920 127130 66972
rect 154482 66920 154488 66972
rect 154540 66960 154546 66972
rect 355226 66960 355232 66972
rect 154540 66932 355232 66960
rect 154540 66920 154546 66932
rect 355226 66920 355232 66932
rect 355284 66920 355290 66972
rect 60826 66852 60832 66904
rect 60884 66892 60890 66904
rect 124398 66892 124404 66904
rect 60884 66864 124404 66892
rect 60884 66852 60890 66864
rect 124398 66852 124404 66864
rect 124456 66852 124462 66904
rect 141694 66852 141700 66904
rect 141752 66892 141758 66904
rect 141878 66892 141884 66904
rect 141752 66864 141884 66892
rect 141752 66852 141758 66864
rect 141878 66852 141884 66864
rect 141936 66852 141942 66904
rect 145558 66852 145564 66904
rect 145616 66892 145622 66904
rect 145926 66892 145932 66904
rect 145616 66864 145932 66892
rect 145616 66852 145622 66864
rect 145926 66852 145932 66864
rect 145984 66852 145990 66904
rect 152182 66852 152188 66904
rect 152240 66892 152246 66904
rect 369394 66892 369400 66904
rect 152240 66864 369400 66892
rect 152240 66852 152246 66864
rect 369394 66852 369400 66864
rect 369452 66852 369458 66904
rect 137094 66716 137100 66768
rect 137152 66756 137158 66768
rect 137738 66756 137744 66768
rect 137152 66728 137744 66756
rect 137152 66716 137158 66728
rect 137738 66716 137744 66728
rect 137796 66716 137802 66768
rect 129182 66240 129188 66292
rect 129240 66280 129246 66292
rect 131298 66280 131304 66292
rect 129240 66252 131304 66280
rect 129240 66240 129246 66252
rect 131298 66240 131304 66252
rect 131356 66240 131362 66292
rect 121914 65968 121920 66020
rect 121972 66008 121978 66020
rect 122190 66008 122196 66020
rect 121972 65980 122196 66008
rect 121972 65968 121978 65980
rect 122190 65968 122196 65980
rect 122248 65968 122254 66020
rect 132862 65968 132868 66020
rect 132920 66008 132926 66020
rect 134610 66008 134616 66020
rect 132920 65980 134616 66008
rect 132920 65968 132926 65980
rect 134610 65968 134616 65980
rect 134668 65968 134674 66020
rect 121546 65900 121552 65952
rect 121604 65940 121610 65952
rect 128262 65940 128268 65952
rect 121604 65912 128268 65940
rect 121604 65900 121610 65912
rect 128262 65900 128268 65912
rect 128320 65900 128326 65952
rect 128814 65900 128820 65952
rect 128872 65940 128878 65952
rect 128998 65940 129004 65952
rect 128872 65912 129004 65940
rect 128872 65900 128878 65912
rect 128998 65900 129004 65912
rect 129056 65900 129062 65952
rect 138750 65900 138756 65952
rect 138808 65940 138814 65952
rect 139210 65940 139216 65952
rect 138808 65912 139216 65940
rect 138808 65900 138814 65912
rect 139210 65900 139216 65912
rect 139268 65900 139274 65952
rect 142706 65900 142712 65952
rect 142764 65940 142770 65952
rect 142982 65940 142988 65952
rect 142764 65912 142988 65940
rect 142764 65900 142770 65912
rect 142982 65900 142988 65912
rect 143040 65900 143046 65952
rect 112438 65832 112444 65884
rect 112496 65872 112502 65884
rect 129918 65872 129924 65884
rect 112496 65844 129924 65872
rect 112496 65832 112502 65844
rect 129918 65832 129924 65844
rect 129976 65832 129982 65884
rect 139946 65832 139952 65884
rect 140004 65872 140010 65884
rect 140406 65872 140412 65884
rect 140004 65844 140412 65872
rect 140004 65832 140010 65844
rect 140406 65832 140412 65844
rect 140464 65832 140470 65884
rect 154942 65832 154948 65884
rect 155000 65872 155006 65884
rect 155770 65872 155776 65884
rect 155000 65844 155776 65872
rect 155000 65832 155006 65844
rect 155770 65832 155776 65844
rect 155828 65832 155834 65884
rect 159726 65832 159732 65884
rect 159784 65872 159790 65884
rect 166902 65872 166908 65884
rect 159784 65844 166908 65872
rect 159784 65832 159790 65844
rect 166902 65832 166908 65844
rect 166960 65832 166966 65884
rect 101030 65764 101036 65816
rect 101088 65804 101094 65816
rect 129366 65804 129372 65816
rect 101088 65776 129372 65804
rect 101088 65764 101094 65776
rect 129366 65764 129372 65776
rect 129424 65764 129430 65816
rect 134242 65764 134248 65816
rect 134300 65804 134306 65816
rect 134886 65804 134892 65816
rect 134300 65776 134892 65804
rect 134300 65764 134306 65776
rect 134886 65764 134892 65776
rect 134944 65764 134950 65816
rect 135070 65764 135076 65816
rect 135128 65804 135134 65816
rect 168374 65804 168380 65816
rect 135128 65776 168380 65804
rect 135128 65764 135134 65776
rect 168374 65764 168380 65776
rect 168432 65764 168438 65816
rect 86862 65696 86868 65748
rect 86920 65736 86926 65748
rect 121546 65736 121552 65748
rect 86920 65708 121552 65736
rect 86920 65696 86926 65708
rect 121546 65696 121552 65708
rect 121604 65696 121610 65748
rect 127894 65736 127900 65748
rect 121748 65708 127900 65736
rect 79686 65628 79692 65680
rect 79744 65668 79750 65680
rect 121748 65668 121776 65708
rect 127894 65696 127900 65708
rect 127952 65696 127958 65748
rect 133414 65736 133420 65748
rect 132604 65708 133420 65736
rect 79744 65640 121776 65668
rect 79744 65628 79750 65640
rect 121822 65628 121828 65680
rect 121880 65668 121886 65680
rect 122374 65668 122380 65680
rect 121880 65640 122380 65668
rect 121880 65628 121886 65640
rect 122374 65628 122380 65640
rect 122432 65628 122438 65680
rect 123294 65628 123300 65680
rect 123352 65668 123358 65680
rect 123938 65668 123944 65680
rect 123352 65640 123944 65668
rect 123352 65628 123358 65640
rect 123938 65628 123944 65640
rect 123996 65628 124002 65680
rect 127526 65628 127532 65680
rect 127584 65668 127590 65680
rect 127802 65668 127808 65680
rect 127584 65640 127808 65668
rect 127584 65628 127590 65640
rect 127802 65628 127808 65640
rect 127860 65628 127866 65680
rect 26510 65560 26516 65612
rect 26568 65600 26574 65612
rect 123110 65600 123116 65612
rect 26568 65572 123116 65600
rect 26568 65560 26574 65572
rect 123110 65560 123116 65572
rect 123168 65560 123174 65612
rect 2866 65492 2872 65544
rect 2924 65532 2930 65544
rect 121638 65532 121644 65544
rect 2924 65504 121644 65532
rect 2924 65492 2930 65504
rect 121638 65492 121644 65504
rect 121696 65492 121702 65544
rect 121730 65492 121736 65544
rect 121788 65532 121794 65544
rect 122558 65532 122564 65544
rect 121788 65504 122564 65532
rect 121788 65492 121794 65504
rect 122558 65492 122564 65504
rect 122616 65492 122622 65544
rect 125134 65492 125140 65544
rect 125192 65532 125198 65544
rect 125502 65532 125508 65544
rect 125192 65504 125508 65532
rect 125192 65492 125198 65504
rect 125502 65492 125508 65504
rect 125560 65492 125566 65544
rect 126146 65492 126152 65544
rect 126204 65532 126210 65544
rect 126606 65532 126612 65544
rect 126204 65504 126612 65532
rect 126204 65492 126210 65504
rect 126606 65492 126612 65504
rect 126664 65492 126670 65544
rect 128722 65492 128728 65544
rect 128780 65532 128786 65544
rect 129274 65532 129280 65544
rect 128780 65504 129280 65532
rect 128780 65492 128786 65504
rect 129274 65492 129280 65504
rect 129332 65492 129338 65544
rect 130654 65492 130660 65544
rect 130712 65532 130718 65544
rect 131574 65532 131580 65544
rect 130712 65504 131580 65532
rect 130712 65492 130718 65504
rect 131574 65492 131580 65504
rect 131632 65492 131638 65544
rect 131942 65492 131948 65544
rect 132000 65532 132006 65544
rect 132310 65532 132316 65544
rect 132000 65504 132316 65532
rect 132000 65492 132006 65504
rect 132310 65492 132316 65504
rect 132368 65492 132374 65544
rect 132604 65408 132632 65708
rect 133414 65696 133420 65708
rect 133472 65696 133478 65748
rect 134334 65696 134340 65748
rect 134392 65736 134398 65748
rect 134794 65736 134800 65748
rect 134392 65708 134800 65736
rect 134392 65696 134398 65708
rect 134794 65696 134800 65708
rect 134852 65696 134858 65748
rect 137094 65696 137100 65748
rect 137152 65736 137158 65748
rect 137646 65736 137652 65748
rect 137152 65708 137652 65736
rect 137152 65696 137158 65708
rect 137646 65696 137652 65708
rect 137704 65696 137710 65748
rect 139762 65696 139768 65748
rect 139820 65736 139826 65748
rect 140314 65736 140320 65748
rect 139820 65708 140320 65736
rect 139820 65696 139826 65708
rect 140314 65696 140320 65708
rect 140372 65696 140378 65748
rect 184198 65736 184204 65748
rect 140424 65708 184204 65736
rect 136818 65628 136824 65680
rect 136876 65668 136882 65680
rect 137462 65668 137468 65680
rect 136876 65640 137468 65668
rect 136876 65628 136882 65640
rect 137462 65628 137468 65640
rect 137520 65628 137526 65680
rect 138382 65628 138388 65680
rect 138440 65628 138446 65680
rect 138566 65628 138572 65680
rect 138624 65628 138630 65680
rect 139394 65628 139400 65680
rect 139452 65668 139458 65680
rect 140424 65668 140452 65708
rect 184198 65696 184204 65708
rect 184256 65696 184262 65748
rect 139452 65640 140452 65668
rect 139452 65628 139458 65640
rect 143994 65628 144000 65680
rect 144052 65668 144058 65680
rect 144270 65668 144276 65680
rect 144052 65640 144276 65668
rect 144052 65628 144058 65640
rect 144270 65628 144276 65640
rect 144328 65628 144334 65680
rect 149330 65628 149336 65680
rect 149388 65668 149394 65680
rect 150158 65668 150164 65680
rect 149388 65640 150164 65668
rect 149388 65628 149394 65640
rect 150158 65628 150164 65640
rect 150216 65628 150222 65680
rect 150526 65628 150532 65680
rect 150584 65668 150590 65680
rect 151262 65668 151268 65680
rect 150584 65640 151268 65668
rect 150584 65628 150590 65640
rect 151262 65628 151268 65640
rect 151320 65628 151326 65680
rect 153562 65628 153568 65680
rect 153620 65668 153626 65680
rect 154390 65668 154396 65680
rect 153620 65640 154396 65668
rect 153620 65628 153626 65640
rect 154390 65628 154396 65640
rect 154448 65628 154454 65680
rect 155126 65628 155132 65680
rect 155184 65668 155190 65680
rect 155184 65640 155448 65668
rect 155184 65628 155190 65640
rect 132770 65600 132776 65612
rect 132696 65572 132776 65600
rect 123478 65356 123484 65408
rect 123536 65396 123542 65408
rect 123846 65396 123852 65408
rect 123536 65368 123852 65396
rect 123536 65356 123542 65368
rect 123846 65356 123852 65368
rect 123904 65356 123910 65408
rect 128998 65356 129004 65408
rect 129056 65396 129062 65408
rect 129182 65396 129188 65408
rect 129056 65368 129188 65396
rect 129056 65356 129062 65368
rect 129182 65356 129188 65368
rect 129240 65356 129246 65408
rect 131850 65356 131856 65408
rect 131908 65396 131914 65408
rect 132126 65396 132132 65408
rect 131908 65368 132132 65396
rect 131908 65356 131914 65368
rect 132126 65356 132132 65368
rect 132184 65356 132190 65408
rect 132586 65356 132592 65408
rect 132644 65356 132650 65408
rect 131758 65288 131764 65340
rect 131816 65288 131822 65340
rect 131776 65136 131804 65288
rect 132696 65260 132724 65572
rect 132770 65560 132776 65572
rect 132828 65560 132834 65612
rect 134058 65560 134064 65612
rect 134116 65600 134122 65612
rect 134426 65600 134432 65612
rect 134116 65572 134432 65600
rect 134116 65560 134122 65572
rect 134426 65560 134432 65572
rect 134484 65560 134490 65612
rect 135622 65560 135628 65612
rect 135680 65600 135686 65612
rect 136174 65600 136180 65612
rect 135680 65572 136180 65600
rect 135680 65560 135686 65572
rect 136174 65560 136180 65572
rect 136232 65560 136238 65612
rect 137278 65560 137284 65612
rect 137336 65600 137342 65612
rect 137646 65600 137652 65612
rect 137336 65572 137652 65600
rect 137336 65560 137342 65572
rect 137646 65560 137652 65572
rect 137704 65560 137710 65612
rect 133966 65492 133972 65544
rect 134024 65532 134030 65544
rect 134978 65532 134984 65544
rect 134024 65504 134984 65532
rect 134024 65492 134030 65504
rect 134978 65492 134984 65504
rect 135036 65492 135042 65544
rect 136910 65492 136916 65544
rect 136968 65532 136974 65544
rect 137462 65532 137468 65544
rect 136968 65504 137468 65532
rect 136968 65492 136974 65504
rect 137462 65492 137468 65504
rect 137520 65492 137526 65544
rect 132770 65356 132776 65408
rect 132828 65396 132834 65408
rect 133414 65396 133420 65408
rect 132828 65368 133420 65396
rect 132828 65356 132834 65368
rect 133414 65356 133420 65368
rect 133472 65356 133478 65408
rect 135346 65356 135352 65408
rect 135404 65396 135410 65408
rect 136082 65396 136088 65408
rect 135404 65368 136088 65396
rect 135404 65356 135410 65368
rect 136082 65356 136088 65368
rect 136140 65356 136146 65408
rect 133414 65260 133420 65272
rect 132696 65232 133420 65260
rect 133414 65220 133420 65232
rect 133472 65220 133478 65272
rect 138400 65192 138428 65628
rect 138584 65396 138612 65628
rect 142246 65560 142252 65612
rect 142304 65600 142310 65612
rect 143258 65600 143264 65612
rect 142304 65572 143264 65600
rect 142304 65560 142310 65572
rect 143258 65560 143264 65572
rect 143316 65560 143322 65612
rect 143626 65560 143632 65612
rect 143684 65600 143690 65612
rect 144546 65600 144552 65612
rect 143684 65572 144552 65600
rect 143684 65560 143690 65572
rect 144546 65560 144552 65572
rect 144604 65560 144610 65612
rect 144914 65560 144920 65612
rect 144972 65600 144978 65612
rect 145742 65600 145748 65612
rect 144972 65572 145748 65600
rect 144972 65560 144978 65572
rect 145742 65560 145748 65572
rect 145800 65560 145806 65612
rect 148042 65560 148048 65612
rect 148100 65600 148106 65612
rect 148778 65600 148784 65612
rect 148100 65572 148784 65600
rect 148100 65560 148106 65572
rect 148778 65560 148784 65572
rect 148836 65560 148842 65612
rect 149882 65600 149888 65612
rect 149440 65572 149888 65600
rect 138934 65492 138940 65544
rect 138992 65532 138998 65544
rect 139118 65532 139124 65544
rect 138992 65504 139124 65532
rect 138992 65492 138998 65504
rect 139118 65492 139124 65504
rect 139176 65492 139182 65544
rect 139486 65492 139492 65544
rect 139544 65532 139550 65544
rect 140498 65532 140504 65544
rect 139544 65504 140504 65532
rect 139544 65492 139550 65504
rect 140498 65492 140504 65504
rect 140556 65492 140562 65544
rect 140866 65492 140872 65544
rect 140924 65532 140930 65544
rect 141786 65532 141792 65544
rect 140924 65504 141792 65532
rect 140924 65492 140930 65504
rect 141786 65492 141792 65504
rect 141844 65492 141850 65544
rect 142430 65492 142436 65544
rect 142488 65532 142494 65544
rect 143166 65532 143172 65544
rect 142488 65504 143172 65532
rect 142488 65492 142494 65504
rect 143166 65492 143172 65504
rect 143224 65492 143230 65544
rect 144086 65492 144092 65544
rect 144144 65532 144150 65544
rect 144638 65532 144644 65544
rect 144144 65504 144644 65532
rect 144144 65492 144150 65504
rect 144638 65492 144644 65504
rect 144696 65492 144702 65544
rect 145190 65492 145196 65544
rect 145248 65532 145254 65544
rect 145834 65532 145840 65544
rect 145248 65504 145840 65532
rect 145248 65492 145254 65504
rect 145834 65492 145840 65504
rect 145892 65492 145898 65544
rect 147674 65492 147680 65544
rect 147732 65532 147738 65544
rect 148134 65532 148140 65544
rect 147732 65504 148140 65532
rect 147732 65492 147738 65504
rect 148134 65492 148140 65504
rect 148192 65492 148198 65544
rect 148318 65492 148324 65544
rect 148376 65532 148382 65544
rect 148686 65532 148692 65544
rect 148376 65504 148692 65532
rect 148376 65492 148382 65504
rect 148686 65492 148692 65504
rect 148744 65492 148750 65544
rect 139854 65424 139860 65476
rect 139912 65464 139918 65476
rect 140222 65464 140228 65476
rect 139912 65436 140228 65464
rect 139912 65424 139918 65436
rect 140222 65424 140228 65436
rect 140280 65424 140286 65476
rect 149440 65408 149468 65572
rect 149882 65560 149888 65572
rect 149940 65560 149946 65612
rect 153194 65560 153200 65612
rect 153252 65600 153258 65612
rect 154022 65600 154028 65612
rect 153252 65572 154028 65600
rect 153252 65560 153258 65572
rect 154022 65560 154028 65572
rect 154080 65560 154086 65612
rect 154666 65560 154672 65612
rect 154724 65600 154730 65612
rect 155218 65600 155224 65612
rect 154724 65572 155224 65600
rect 154724 65560 154730 65572
rect 155218 65560 155224 65572
rect 155276 65560 155282 65612
rect 149606 65492 149612 65544
rect 149664 65532 149670 65544
rect 149974 65532 149980 65544
rect 149664 65504 149980 65532
rect 149664 65492 149670 65504
rect 149974 65492 149980 65504
rect 150032 65492 150038 65544
rect 150526 65492 150532 65544
rect 150584 65532 150590 65544
rect 150986 65532 150992 65544
rect 150584 65504 150992 65532
rect 150584 65492 150590 65504
rect 150986 65492 150992 65504
rect 151044 65492 151050 65544
rect 151814 65492 151820 65544
rect 151872 65532 151878 65544
rect 152918 65532 152924 65544
rect 151872 65504 152924 65532
rect 151872 65492 151878 65504
rect 152918 65492 152924 65504
rect 152976 65492 152982 65544
rect 153746 65492 153752 65544
rect 153804 65532 153810 65544
rect 154206 65532 154212 65544
rect 153804 65504 154212 65532
rect 153804 65492 153810 65504
rect 154206 65492 154212 65504
rect 154264 65492 154270 65544
rect 151170 65464 151176 65476
rect 151096 65436 151176 65464
rect 138934 65396 138940 65408
rect 138584 65368 138940 65396
rect 138934 65356 138940 65368
rect 138992 65356 138998 65408
rect 143902 65356 143908 65408
rect 143960 65396 143966 65408
rect 144362 65396 144368 65408
rect 143960 65368 144368 65396
rect 143960 65356 143966 65368
rect 144362 65356 144368 65368
rect 144420 65356 144426 65408
rect 146662 65356 146668 65408
rect 146720 65396 146726 65408
rect 147214 65396 147220 65408
rect 146720 65368 147220 65396
rect 146720 65356 146726 65368
rect 147214 65356 147220 65368
rect 147272 65356 147278 65408
rect 149422 65356 149428 65408
rect 149480 65356 149486 65408
rect 146846 65288 146852 65340
rect 146904 65328 146910 65340
rect 147306 65328 147312 65340
rect 146904 65300 147312 65328
rect 146904 65288 146910 65300
rect 147306 65288 147312 65300
rect 147364 65288 147370 65340
rect 151096 65272 151124 65436
rect 151170 65424 151176 65436
rect 151228 65424 151234 65476
rect 153470 65424 153476 65476
rect 153528 65464 153534 65476
rect 154298 65464 154304 65476
rect 153528 65436 154304 65464
rect 153528 65424 153534 65436
rect 154298 65424 154304 65436
rect 154356 65424 154362 65476
rect 155420 65408 155448 65640
rect 156230 65628 156236 65680
rect 156288 65668 156294 65680
rect 446214 65668 446220 65680
rect 156288 65640 446220 65668
rect 156288 65628 156294 65640
rect 446214 65628 446220 65640
rect 446272 65628 446278 65680
rect 160094 65560 160100 65612
rect 160152 65600 160158 65612
rect 161106 65600 161112 65612
rect 160152 65572 161112 65600
rect 160152 65560 160158 65572
rect 161106 65560 161112 65572
rect 161164 65560 161170 65612
rect 162026 65560 162032 65612
rect 162084 65600 162090 65612
rect 162486 65600 162492 65612
rect 162084 65572 162492 65600
rect 162084 65560 162090 65572
rect 162486 65560 162492 65572
rect 162544 65560 162550 65612
rect 163222 65560 163228 65612
rect 163280 65600 163286 65612
rect 163682 65600 163688 65612
rect 163280 65572 163688 65600
rect 163280 65560 163286 65572
rect 163682 65560 163688 65572
rect 163740 65560 163746 65612
rect 164234 65560 164240 65612
rect 164292 65600 164298 65612
rect 165246 65600 165252 65612
rect 164292 65572 165252 65600
rect 164292 65560 164298 65572
rect 165246 65560 165252 65572
rect 165304 65560 165310 65612
rect 165614 65560 165620 65612
rect 165672 65600 165678 65612
rect 166718 65600 166724 65612
rect 165672 65572 166724 65600
rect 165672 65560 165678 65572
rect 166718 65560 166724 65572
rect 166776 65560 166782 65612
rect 487614 65600 487620 65612
rect 166828 65572 487620 65600
rect 157426 65492 157432 65544
rect 157484 65532 157490 65544
rect 157886 65532 157892 65544
rect 157484 65504 157892 65532
rect 157484 65492 157490 65504
rect 157886 65492 157892 65504
rect 157944 65492 157950 65544
rect 158714 65492 158720 65544
rect 158772 65532 158778 65544
rect 159174 65532 159180 65544
rect 158772 65504 159180 65532
rect 158772 65492 158778 65504
rect 159174 65492 159180 65504
rect 159232 65492 159238 65544
rect 160462 65492 160468 65544
rect 160520 65532 160526 65544
rect 160830 65532 160836 65544
rect 160520 65504 160836 65532
rect 160520 65492 160526 65504
rect 160830 65492 160836 65504
rect 160888 65492 160894 65544
rect 162854 65492 162860 65544
rect 162912 65532 162918 65544
rect 164050 65532 164056 65544
rect 162912 65504 164056 65532
rect 162912 65492 162918 65504
rect 164050 65492 164056 65504
rect 164108 65492 164114 65544
rect 164510 65492 164516 65544
rect 164568 65532 164574 65544
rect 165062 65532 165068 65544
rect 164568 65504 165068 65532
rect 164568 65492 164574 65504
rect 165062 65492 165068 65504
rect 165120 65492 165126 65544
rect 165798 65492 165804 65544
rect 165856 65532 165862 65544
rect 166534 65532 166540 65544
rect 165856 65504 166540 65532
rect 165856 65492 165862 65504
rect 166534 65492 166540 65504
rect 166592 65492 166598 65544
rect 160002 65424 160008 65476
rect 160060 65464 160066 65476
rect 160060 65436 164004 65464
rect 160060 65424 160066 65436
rect 155402 65356 155408 65408
rect 155460 65356 155466 65408
rect 159266 65356 159272 65408
rect 159324 65396 159330 65408
rect 159726 65396 159732 65408
rect 159324 65368 159732 65396
rect 159324 65356 159330 65368
rect 159726 65356 159732 65368
rect 159784 65356 159790 65408
rect 163406 65356 163412 65408
rect 163464 65396 163470 65408
rect 163866 65396 163872 65408
rect 163464 65368 163872 65396
rect 163464 65356 163470 65368
rect 163866 65356 163872 65368
rect 163924 65356 163930 65408
rect 163976 65396 164004 65436
rect 164326 65424 164332 65476
rect 164384 65464 164390 65476
rect 165338 65464 165344 65476
rect 164384 65436 165344 65464
rect 164384 65424 164390 65436
rect 165338 65424 165344 65436
rect 165396 65424 165402 65476
rect 166828 65464 166856 65572
rect 487614 65560 487620 65572
rect 487672 65560 487678 65612
rect 166902 65492 166908 65544
rect 166960 65532 166966 65544
rect 491110 65532 491116 65544
rect 166960 65504 491116 65532
rect 166960 65492 166966 65504
rect 491110 65492 491116 65504
rect 491168 65492 491174 65544
rect 165448 65436 166856 65464
rect 165448 65396 165476 65436
rect 163976 65368 165476 65396
rect 165706 65356 165712 65408
rect 165764 65396 165770 65408
rect 166258 65396 166264 65408
rect 165764 65368 166264 65396
rect 165764 65356 165770 65368
rect 166258 65356 166264 65368
rect 166316 65356 166322 65408
rect 154850 65288 154856 65340
rect 154908 65328 154914 65340
rect 155586 65328 155592 65340
rect 154908 65300 155592 65328
rect 154908 65288 154914 65300
rect 155586 65288 155592 65300
rect 155644 65288 155650 65340
rect 163314 65288 163320 65340
rect 163372 65328 163378 65340
rect 163774 65328 163780 65340
rect 163372 65300 163780 65328
rect 163372 65288 163378 65300
rect 163774 65288 163780 65300
rect 163832 65288 163838 65340
rect 138658 65220 138664 65272
rect 138716 65260 138722 65272
rect 139026 65260 139032 65272
rect 138716 65232 139032 65260
rect 138716 65220 138722 65232
rect 139026 65220 139032 65232
rect 139084 65220 139090 65272
rect 139578 65220 139584 65272
rect 139636 65260 139642 65272
rect 140314 65260 140320 65272
rect 139636 65232 140320 65260
rect 139636 65220 139642 65232
rect 140314 65220 140320 65232
rect 140372 65220 140378 65272
rect 142522 65220 142528 65272
rect 142580 65260 142586 65272
rect 142890 65260 142896 65272
rect 142580 65232 142896 65260
rect 142580 65220 142586 65232
rect 142890 65220 142896 65232
rect 142948 65220 142954 65272
rect 146294 65220 146300 65272
rect 146352 65260 146358 65272
rect 147122 65260 147128 65272
rect 146352 65232 147128 65260
rect 146352 65220 146358 65232
rect 147122 65220 147128 65232
rect 147180 65220 147186 65272
rect 147858 65220 147864 65272
rect 147916 65260 147922 65272
rect 148318 65260 148324 65272
rect 147916 65232 148324 65260
rect 147916 65220 147922 65232
rect 148318 65220 148324 65232
rect 148376 65220 148382 65272
rect 151078 65220 151084 65272
rect 151136 65220 151142 65272
rect 154574 65220 154580 65272
rect 154632 65260 154638 65272
rect 155494 65260 155500 65272
rect 154632 65232 155500 65260
rect 154632 65220 154638 65232
rect 155494 65220 155500 65232
rect 155552 65220 155558 65272
rect 158898 65220 158904 65272
rect 158956 65260 158962 65272
rect 159358 65260 159364 65272
rect 158956 65232 159364 65260
rect 158956 65220 158962 65232
rect 159358 65220 159364 65232
rect 159416 65220 159422 65272
rect 161658 65220 161664 65272
rect 161716 65260 161722 65272
rect 162210 65260 162216 65272
rect 161716 65232 162216 65260
rect 161716 65220 161722 65232
rect 162210 65220 162216 65232
rect 162268 65220 162274 65272
rect 162946 65220 162952 65272
rect 163004 65260 163010 65272
rect 163866 65260 163872 65272
rect 163004 65232 163872 65260
rect 163004 65220 163010 65232
rect 163866 65220 163872 65232
rect 163924 65220 163930 65272
rect 138750 65192 138756 65204
rect 138400 65164 138756 65192
rect 138750 65152 138756 65164
rect 138808 65152 138814 65204
rect 158990 65152 158996 65204
rect 159048 65192 159054 65204
rect 159542 65192 159548 65204
rect 159048 65164 159548 65192
rect 159048 65152 159054 65164
rect 159542 65152 159548 65164
rect 159600 65152 159606 65204
rect 131758 65084 131764 65136
rect 131816 65084 131822 65136
rect 138014 65084 138020 65136
rect 138072 65124 138078 65136
rect 138842 65124 138848 65136
rect 138072 65096 138848 65124
rect 138072 65084 138078 65096
rect 138842 65084 138848 65096
rect 138900 65084 138906 65136
rect 158806 65084 158812 65136
rect 158864 65124 158870 65136
rect 159450 65124 159456 65136
rect 158864 65096 159456 65124
rect 158864 65084 158870 65096
rect 159450 65084 159456 65096
rect 159508 65084 159514 65136
rect 138198 64948 138204 65000
rect 138256 64988 138262 65000
rect 138934 64988 138940 65000
rect 138256 64960 138940 64988
rect 138256 64948 138262 64960
rect 138934 64948 138940 64960
rect 138992 64948 138998 65000
rect 112806 64336 112812 64388
rect 112864 64376 112870 64388
rect 130562 64376 130568 64388
rect 112864 64348 130568 64376
rect 112864 64336 112870 64348
rect 130562 64336 130568 64348
rect 130620 64336 130626 64388
rect 67910 64268 67916 64320
rect 67968 64308 67974 64320
rect 124122 64308 124128 64320
rect 67968 64280 124128 64308
rect 67968 64268 67974 64280
rect 124122 64268 124128 64280
rect 124180 64268 124186 64320
rect 135714 64268 135720 64320
rect 135772 64308 135778 64320
rect 178678 64308 178684 64320
rect 135772 64280 178684 64308
rect 135772 64268 135778 64280
rect 178678 64268 178684 64280
rect 178736 64268 178742 64320
rect 48958 64200 48964 64252
rect 49016 64240 49022 64252
rect 125318 64240 125324 64252
rect 49016 64212 125324 64240
rect 49016 64200 49022 64212
rect 125318 64200 125324 64212
rect 125376 64200 125382 64252
rect 152366 64200 152372 64252
rect 152424 64200 152430 64252
rect 152458 64200 152464 64252
rect 152516 64240 152522 64252
rect 397730 64240 397736 64252
rect 152516 64212 397736 64240
rect 152516 64200 152522 64212
rect 397730 64200 397736 64212
rect 397788 64200 397794 64252
rect 12342 64132 12348 64184
rect 12400 64172 12406 64184
rect 122466 64172 122472 64184
rect 12400 64144 122472 64172
rect 12400 64132 12406 64144
rect 122466 64132 122472 64144
rect 122524 64132 122530 64184
rect 152384 64048 152412 64200
rect 162670 64132 162676 64184
rect 162728 64172 162734 64184
rect 519538 64172 519544 64184
rect 162728 64144 519544 64172
rect 162728 64132 162734 64144
rect 519538 64132 519544 64144
rect 519596 64132 519602 64184
rect 152366 63996 152372 64048
rect 152424 63996 152430 64048
rect 146386 63724 146392 63776
rect 146444 63764 146450 63776
rect 147030 63764 147036 63776
rect 146444 63736 147036 63764
rect 146444 63724 146450 63736
rect 147030 63724 147036 63736
rect 147088 63724 147094 63776
rect 161842 63452 161848 63504
rect 161900 63492 161906 63504
rect 162394 63492 162400 63504
rect 161900 63464 162400 63492
rect 161900 63452 161906 63464
rect 162394 63452 162400 63464
rect 162452 63452 162458 63504
rect 156414 63316 156420 63368
rect 156472 63356 156478 63368
rect 157058 63356 157064 63368
rect 156472 63328 157064 63356
rect 156472 63316 156478 63328
rect 157058 63316 157064 63328
rect 157116 63316 157122 63368
rect 137738 63044 137744 63096
rect 137796 63084 137802 63096
rect 200298 63084 200304 63096
rect 137796 63056 200304 63084
rect 137796 63044 137802 63056
rect 200298 63044 200304 63056
rect 200356 63044 200362 63096
rect 4798 62976 4804 63028
rect 4856 63016 4862 63028
rect 170306 63016 170312 63028
rect 4856 62988 170312 63016
rect 4856 62976 4862 62988
rect 170306 62976 170312 62988
rect 170364 62976 170370 63028
rect 102226 62908 102232 62960
rect 102284 62948 102290 62960
rect 129458 62948 129464 62960
rect 102284 62920 129464 62948
rect 102284 62908 102290 62920
rect 129458 62908 129464 62920
rect 129516 62908 129522 62960
rect 136726 62908 136732 62960
rect 136784 62948 136790 62960
rect 137738 62948 137744 62960
rect 136784 62920 137744 62948
rect 136784 62908 136790 62920
rect 137738 62908 137744 62920
rect 137796 62908 137802 62960
rect 149054 62908 149060 62960
rect 149112 62948 149118 62960
rect 356330 62948 356336 62960
rect 149112 62920 356336 62948
rect 149112 62908 149118 62920
rect 356330 62908 356336 62920
rect 356388 62908 356394 62960
rect 56042 62840 56048 62892
rect 56100 62880 56106 62892
rect 125870 62880 125876 62892
rect 56100 62852 125876 62880
rect 56100 62840 56106 62852
rect 125870 62840 125876 62852
rect 125928 62840 125934 62892
rect 158254 62840 158260 62892
rect 158312 62880 158318 62892
rect 394234 62880 394240 62892
rect 158312 62852 394240 62880
rect 158312 62840 158318 62852
rect 394234 62840 394240 62852
rect 394292 62840 394298 62892
rect 44266 62772 44272 62824
rect 44324 62812 44330 62824
rect 124950 62812 124956 62824
rect 44324 62784 124956 62812
rect 44324 62772 44330 62784
rect 124950 62772 124956 62784
rect 125008 62772 125014 62824
rect 162762 62772 162768 62824
rect 162820 62812 162826 62824
rect 523034 62812 523040 62824
rect 162820 62784 523040 62812
rect 162820 62772 162826 62784
rect 523034 62772 523040 62784
rect 523092 62772 523098 62824
rect 133230 62024 133236 62076
rect 133288 62064 133294 62076
rect 135990 62064 135996 62076
rect 133288 62036 135996 62064
rect 133288 62024 133294 62036
rect 135990 62024 135996 62036
rect 136048 62024 136054 62076
rect 109310 61480 109316 61532
rect 109368 61520 109374 61532
rect 130010 61520 130016 61532
rect 109368 61492 130016 61520
rect 109368 61480 109374 61492
rect 130010 61480 130016 61492
rect 130068 61480 130074 61532
rect 139210 61480 139216 61532
rect 139268 61520 139274 61532
rect 221550 61520 221556 61532
rect 139268 61492 221556 61520
rect 139268 61480 139274 61492
rect 221550 61480 221556 61492
rect 221608 61480 221614 61532
rect 65518 61412 65524 61464
rect 65576 61452 65582 61464
rect 126698 61452 126704 61464
rect 65576 61424 126704 61452
rect 65576 61412 65582 61424
rect 126698 61412 126704 61424
rect 126756 61412 126762 61464
rect 150618 61412 150624 61464
rect 150676 61452 150682 61464
rect 374086 61452 374092 61464
rect 150676 61424 374092 61452
rect 150676 61412 150682 61424
rect 374086 61412 374092 61424
rect 374144 61412 374150 61464
rect 40678 61344 40684 61396
rect 40736 61384 40742 61396
rect 124674 61384 124680 61396
rect 40736 61356 124680 61384
rect 40736 61344 40742 61356
rect 124674 61344 124680 61356
rect 124732 61344 124738 61396
rect 156690 61344 156696 61396
rect 156748 61384 156754 61396
rect 453298 61384 453304 61396
rect 156748 61356 453304 61384
rect 156748 61344 156754 61356
rect 453298 61344 453304 61356
rect 453356 61344 453362 61396
rect 157702 61140 157708 61192
rect 157760 61180 157766 61192
rect 157978 61180 157984 61192
rect 157760 61152 157984 61180
rect 157760 61140 157766 61152
rect 157978 61140 157984 61152
rect 158036 61140 158042 61192
rect 149790 61072 149796 61124
rect 149848 61112 149854 61124
rect 150066 61112 150072 61124
rect 149848 61084 150072 61112
rect 149848 61072 149854 61084
rect 150066 61072 150072 61084
rect 150124 61072 150130 61124
rect 117222 60800 117228 60852
rect 117280 60840 117286 60852
rect 122282 60840 122288 60852
rect 117280 60812 122288 60840
rect 117280 60800 117286 60812
rect 122282 60800 122288 60812
rect 122340 60800 122346 60852
rect 137186 60188 137192 60240
rect 137244 60228 137250 60240
rect 207382 60228 207388 60240
rect 137244 60200 207388 60228
rect 137244 60188 137250 60200
rect 207382 60188 207388 60200
rect 207440 60188 207446 60240
rect 63218 60120 63224 60172
rect 63276 60160 63282 60172
rect 126790 60160 126796 60172
rect 63276 60132 126796 60160
rect 63276 60120 63282 60132
rect 126790 60120 126796 60132
rect 126848 60120 126854 60172
rect 140130 60120 140136 60172
rect 140188 60160 140194 60172
rect 239306 60160 239312 60172
rect 140188 60132 239312 60160
rect 140188 60120 140194 60132
rect 239306 60120 239312 60132
rect 239364 60120 239370 60172
rect 59630 60052 59636 60104
rect 59688 60092 59694 60104
rect 126606 60092 126612 60104
rect 59688 60064 126612 60092
rect 59688 60052 59694 60064
rect 126606 60052 126612 60064
rect 126664 60052 126670 60104
rect 148318 60052 148324 60104
rect 148376 60092 148382 60104
rect 338666 60092 338672 60104
rect 148376 60064 338672 60092
rect 148376 60052 148382 60064
rect 338666 60052 338672 60064
rect 338724 60052 338730 60104
rect 9950 59984 9956 60036
rect 10008 60024 10014 60036
rect 117222 60024 117228 60036
rect 10008 59996 117228 60024
rect 10008 59984 10014 59996
rect 117222 59984 117228 59996
rect 117280 59984 117286 60036
rect 126238 59984 126244 60036
rect 126296 60024 126302 60036
rect 130838 60024 130844 60036
rect 126296 59996 130844 60024
rect 126296 59984 126302 59996
rect 130838 59984 130844 59996
rect 130896 59984 130902 60036
rect 151078 59984 151084 60036
rect 151136 60024 151142 60036
rect 381170 60024 381176 60036
rect 151136 59996 381176 60024
rect 151136 59984 151142 59996
rect 381170 59984 381176 59996
rect 381228 59984 381234 60036
rect 135254 58896 135260 58948
rect 135312 58936 135318 58948
rect 176654 58936 176660 58948
rect 135312 58908 176660 58936
rect 135312 58896 135318 58908
rect 176654 58896 176660 58908
rect 176712 58896 176718 58948
rect 152458 58828 152464 58880
rect 152516 58868 152522 58880
rect 277118 58868 277124 58880
rect 152516 58840 277124 58868
rect 152516 58828 152522 58840
rect 277118 58828 277124 58840
rect 277176 58828 277182 58880
rect 153930 58760 153936 58812
rect 153988 58800 153994 58812
rect 409598 58800 409604 58812
rect 153988 58772 409604 58800
rect 153988 58760 153994 58772
rect 409598 58760 409604 58772
rect 409656 58760 409662 58812
rect 163406 58692 163412 58744
rect 163464 58732 163470 58744
rect 544378 58732 544384 58744
rect 163464 58704 544384 58732
rect 163464 58692 163470 58704
rect 544378 58692 544384 58704
rect 544436 58692 544442 58744
rect 25314 58624 25320 58676
rect 25372 58664 25378 58676
rect 123846 58664 123852 58676
rect 25372 58636 123852 58664
rect 25372 58624 25378 58636
rect 123846 58624 123852 58636
rect 123904 58624 123910 58676
rect 166442 58624 166448 58676
rect 166500 58664 166506 58676
rect 572714 58664 572720 58676
rect 166500 58636 572720 58664
rect 166500 58624 166506 58636
rect 572714 58624 572720 58636
rect 572772 58624 572778 58676
rect 114002 58352 114008 58404
rect 114060 58392 114066 58404
rect 119614 58392 119620 58404
rect 114060 58364 119620 58392
rect 114060 58352 114066 58364
rect 119614 58352 119620 58364
rect 119672 58352 119678 58404
rect 133230 57876 133236 57928
rect 133288 57916 133294 57928
rect 136358 57916 136364 57928
rect 133288 57888 136364 57916
rect 133288 57876 133294 57888
rect 136358 57876 136364 57888
rect 136416 57876 136422 57928
rect 138658 57400 138664 57452
rect 138716 57440 138722 57452
rect 225138 57440 225144 57452
rect 138716 57412 225144 57440
rect 138716 57400 138722 57412
rect 225138 57400 225144 57412
rect 225196 57400 225202 57452
rect 106918 57332 106924 57384
rect 106976 57372 106982 57384
rect 121270 57372 121276 57384
rect 106976 57344 121276 57372
rect 106976 57332 106982 57344
rect 121270 57332 121276 57344
rect 121328 57332 121334 57384
rect 142706 57332 142712 57384
rect 142764 57372 142770 57384
rect 271230 57372 271236 57384
rect 142764 57344 271236 57372
rect 142764 57332 142770 57344
rect 271230 57332 271236 57344
rect 271288 57332 271294 57384
rect 77386 57264 77392 57316
rect 77444 57304 77450 57316
rect 127802 57304 127808 57316
rect 77444 57276 127808 57304
rect 77444 57264 77450 57276
rect 127802 57264 127808 57276
rect 127860 57264 127866 57316
rect 145558 57264 145564 57316
rect 145616 57304 145622 57316
rect 313826 57304 313832 57316
rect 145616 57276 313832 57304
rect 145616 57264 145622 57276
rect 313826 57264 313832 57276
rect 313884 57264 313890 57316
rect 8754 57196 8760 57248
rect 8812 57236 8818 57248
rect 121822 57236 121828 57248
rect 8812 57208 121828 57236
rect 8812 57196 8818 57208
rect 121822 57196 121828 57208
rect 121880 57196 121886 57248
rect 163498 57196 163504 57248
rect 163556 57236 163562 57248
rect 540790 57236 540796 57248
rect 163556 57208 540796 57236
rect 163556 57196 163562 57208
rect 540790 57196 540796 57208
rect 540848 57196 540854 57248
rect 136082 55972 136088 56024
rect 136140 56012 136146 56024
rect 177850 56012 177856 56024
rect 136140 55984 177856 56012
rect 136140 55972 136146 55984
rect 177850 55972 177856 55984
rect 177908 55972 177914 56024
rect 57238 55904 57244 55956
rect 57296 55944 57302 55956
rect 123570 55944 123576 55956
rect 57296 55916 123576 55944
rect 57296 55904 57302 55916
rect 123570 55904 123576 55916
rect 123628 55904 123634 55956
rect 149606 55904 149612 55956
rect 149664 55944 149670 55956
rect 359918 55944 359924 55956
rect 149664 55916 359924 55944
rect 149664 55904 149670 55916
rect 359918 55904 359924 55916
rect 359976 55904 359982 55956
rect 32398 55836 32404 55888
rect 32456 55876 32462 55888
rect 123754 55876 123760 55888
rect 32456 55848 123760 55876
rect 32456 55836 32462 55848
rect 123754 55836 123760 55848
rect 123812 55836 123818 55888
rect 164970 55836 164976 55888
rect 165028 55876 165034 55888
rect 558546 55876 558552 55888
rect 165028 55848 558552 55876
rect 165028 55836 165034 55848
rect 558546 55836 558552 55848
rect 558604 55836 558610 55888
rect 138750 54748 138756 54800
rect 138808 54788 138814 54800
rect 216858 54788 216864 54800
rect 138808 54760 216864 54788
rect 138808 54748 138814 54760
rect 216858 54748 216864 54760
rect 216916 54748 216922 54800
rect 142798 54680 142804 54732
rect 142856 54720 142862 54732
rect 274818 54720 274824 54732
rect 142856 54692 274824 54720
rect 142856 54680 142862 54692
rect 274818 54680 274824 54692
rect 274876 54680 274882 54732
rect 146846 54612 146852 54664
rect 146904 54652 146910 54664
rect 324406 54652 324412 54664
rect 146904 54624 324412 54652
rect 146904 54612 146910 54624
rect 324406 54612 324412 54624
rect 324464 54612 324470 54664
rect 155126 54544 155132 54596
rect 155184 54584 155190 54596
rect 427262 54584 427268 54596
rect 155184 54556 427268 54584
rect 155184 54544 155190 54556
rect 427262 54544 427268 54556
rect 427320 54544 427326 54596
rect 33594 54476 33600 54528
rect 33652 54516 33658 54528
rect 123386 54516 123392 54528
rect 33652 54488 123392 54516
rect 33652 54476 33658 54488
rect 123386 54476 123392 54488
rect 123444 54476 123450 54528
rect 159450 54476 159456 54528
rect 159508 54516 159514 54528
rect 468662 54516 468668 54528
rect 159508 54488 468668 54516
rect 159508 54476 159514 54488
rect 468662 54476 468668 54488
rect 468720 54476 468726 54528
rect 136174 53456 136180 53508
rect 136232 53496 136238 53508
rect 186130 53496 186136 53508
rect 136232 53468 186136 53496
rect 136232 53456 136238 53468
rect 186130 53456 186136 53468
rect 186188 53456 186194 53508
rect 137278 53388 137284 53440
rect 137336 53428 137342 53440
rect 201494 53428 201500 53440
rect 137336 53400 201500 53428
rect 137336 53388 137342 53400
rect 201494 53388 201500 53400
rect 201552 53388 201558 53440
rect 148410 53320 148416 53372
rect 148468 53360 148474 53372
rect 342162 53360 342168 53372
rect 148468 53332 342168 53360
rect 148468 53320 148474 53332
rect 342162 53320 342168 53332
rect 342220 53320 342226 53372
rect 154022 53252 154028 53304
rect 154080 53292 154086 53304
rect 413094 53292 413100 53304
rect 154080 53264 413100 53292
rect 154080 53252 154086 53264
rect 413094 53252 413100 53264
rect 413152 53252 413158 53304
rect 163590 53184 163596 53236
rect 163648 53224 163654 53236
rect 539594 53224 539600 53236
rect 163648 53196 539600 53224
rect 163648 53184 163654 53196
rect 539594 53184 539600 53196
rect 539652 53184 539658 53236
rect 62022 53116 62028 53168
rect 62080 53156 62086 53168
rect 126330 53156 126336 53168
rect 62080 53128 126336 53156
rect 62080 53116 62086 53128
rect 126330 53116 126336 53128
rect 126388 53116 126394 53168
rect 165062 53116 165068 53168
rect 165120 53156 165126 53168
rect 552658 53156 552664 53168
rect 165120 53128 552664 53156
rect 165120 53116 165126 53128
rect 552658 53116 552664 53128
rect 552716 53116 552722 53168
rect 31294 53048 31300 53100
rect 31352 53088 31358 53100
rect 123294 53088 123300 53100
rect 31352 53060 123300 53088
rect 31352 53048 31358 53060
rect 123294 53048 123300 53060
rect 123352 53048 123358 53100
rect 166534 53048 166540 53100
rect 166592 53088 166598 53100
rect 569126 53088 569132 53100
rect 166592 53060 569132 53088
rect 166592 53048 166598 53060
rect 569126 53048 569132 53060
rect 569184 53048 569190 53100
rect 133322 52436 133328 52488
rect 133380 52476 133386 52488
rect 136174 52476 136180 52488
rect 133380 52448 136180 52476
rect 133380 52436 133386 52448
rect 136174 52436 136180 52448
rect 136232 52436 136238 52488
rect 132034 52368 132040 52420
rect 132092 52408 132098 52420
rect 134702 52408 134708 52420
rect 132092 52380 134708 52408
rect 132092 52368 132098 52380
rect 134702 52368 134708 52380
rect 134760 52368 134766 52420
rect 146938 51892 146944 51944
rect 146996 51932 147002 51944
rect 327994 51932 328000 51944
rect 146996 51904 328000 51932
rect 146996 51892 147002 51904
rect 327994 51892 328000 51904
rect 328052 51892 328058 51944
rect 151170 51824 151176 51876
rect 151228 51864 151234 51876
rect 377674 51864 377680 51876
rect 151228 51836 377680 51864
rect 151228 51824 151234 51836
rect 377674 51824 377680 51836
rect 377732 51824 377738 51876
rect 167546 51756 167552 51808
rect 167604 51796 167610 51808
rect 436738 51796 436744 51808
rect 167604 51768 436744 51796
rect 167604 51756 167610 51768
rect 436738 51756 436744 51768
rect 436796 51756 436802 51808
rect 13538 51688 13544 51740
rect 13596 51728 13602 51740
rect 121730 51728 121736 51740
rect 13596 51700 121736 51728
rect 13596 51688 13602 51700
rect 121730 51688 121736 51700
rect 121788 51688 121794 51740
rect 162118 51688 162124 51740
rect 162176 51728 162182 51740
rect 508498 51728 508504 51740
rect 162176 51700 508504 51728
rect 162176 51688 162182 51700
rect 508498 51688 508504 51700
rect 508556 51688 508562 51740
rect 137370 50600 137376 50652
rect 137428 50640 137434 50652
rect 203886 50640 203892 50652
rect 137428 50612 203892 50640
rect 137428 50600 137434 50612
rect 203886 50600 203892 50612
rect 203944 50600 203950 50652
rect 145650 50532 145656 50584
rect 145708 50572 145714 50584
rect 310238 50572 310244 50584
rect 145708 50544 310244 50572
rect 145708 50532 145714 50544
rect 310238 50532 310244 50544
rect 310296 50532 310302 50584
rect 149790 50464 149796 50516
rect 149848 50504 149854 50516
rect 367002 50504 367008 50516
rect 149848 50476 367008 50504
rect 149848 50464 149854 50476
rect 367002 50464 367008 50476
rect 367060 50464 367066 50516
rect 155218 50396 155224 50448
rect 155276 50436 155282 50448
rect 430850 50436 430856 50448
rect 155276 50408 430856 50436
rect 155276 50396 155282 50408
rect 430850 50396 430856 50408
rect 430908 50396 430914 50448
rect 14734 50328 14740 50380
rect 14792 50368 14798 50380
rect 122650 50368 122656 50380
rect 14792 50340 122656 50368
rect 14792 50328 14798 50340
rect 122650 50328 122656 50340
rect 122708 50328 122714 50380
rect 165154 50328 165160 50380
rect 165212 50368 165218 50380
rect 562042 50368 562048 50380
rect 165212 50340 562048 50368
rect 165212 50328 165218 50340
rect 562042 50328 562048 50340
rect 562100 50328 562106 50380
rect 136266 49036 136272 49088
rect 136324 49076 136330 49088
rect 184934 49076 184940 49088
rect 136324 49048 184940 49076
rect 136324 49036 136330 49048
rect 184934 49036 184940 49048
rect 184992 49036 184998 49088
rect 99834 48968 99840 49020
rect 99892 49008 99898 49020
rect 121178 49008 121184 49020
rect 99892 48980 121184 49008
rect 99892 48968 99898 48980
rect 121178 48968 121184 48980
rect 121236 48968 121242 49020
rect 148502 48968 148508 49020
rect 148560 49008 148566 49020
rect 345750 49008 345756 49020
rect 148560 48980 345756 49008
rect 148560 48968 148566 48980
rect 345750 48968 345756 48980
rect 345808 48968 345814 49020
rect 135438 47812 135444 47864
rect 135496 47852 135502 47864
rect 180242 47852 180248 47864
rect 135496 47824 180248 47852
rect 135496 47812 135502 47824
rect 180242 47812 180248 47824
rect 180300 47812 180306 47864
rect 144178 47744 144184 47796
rect 144236 47784 144242 47796
rect 291378 47784 291384 47796
rect 144236 47756 291384 47784
rect 144236 47744 144242 47756
rect 291378 47744 291384 47756
rect 291436 47744 291442 47796
rect 149882 47676 149888 47728
rect 149940 47716 149946 47728
rect 363506 47716 363512 47728
rect 149940 47688 363512 47716
rect 149940 47676 149946 47688
rect 363506 47676 363512 47688
rect 363564 47676 363570 47728
rect 92750 47608 92756 47660
rect 92808 47648 92814 47660
rect 129274 47648 129280 47660
rect 92808 47620 129280 47648
rect 92808 47608 92814 47620
rect 129274 47608 129280 47620
rect 129332 47608 129338 47660
rect 154114 47608 154120 47660
rect 154172 47648 154178 47660
rect 416682 47648 416688 47660
rect 154172 47620 416688 47648
rect 154172 47608 154178 47620
rect 416682 47608 416688 47620
rect 416740 47608 416746 47660
rect 83274 47540 83280 47592
rect 83332 47580 83338 47592
rect 127986 47580 127992 47592
rect 83332 47552 127992 47580
rect 83332 47540 83338 47552
rect 127986 47540 127992 47552
rect 128044 47540 128050 47592
rect 156782 47540 156788 47592
rect 156840 47580 156846 47592
rect 442626 47580 442632 47592
rect 156840 47552 442632 47580
rect 156840 47540 156846 47552
rect 442626 47540 442632 47552
rect 442684 47540 442690 47592
rect 135622 46248 135628 46300
rect 135680 46288 135686 46300
rect 188522 46288 188528 46300
rect 135680 46260 188528 46288
rect 135680 46248 135686 46260
rect 188522 46248 188528 46260
rect 188580 46248 188586 46300
rect 4062 46180 4068 46232
rect 4120 46220 4126 46232
rect 122282 46220 122288 46232
rect 4120 46192 122288 46220
rect 4120 46180 4126 46192
rect 122282 46180 122288 46192
rect 122340 46180 122346 46232
rect 140222 46180 140228 46232
rect 140280 46220 140286 46232
rect 234614 46220 234620 46232
rect 140280 46192 234620 46220
rect 140280 46180 140286 46192
rect 234614 46180 234620 46192
rect 234672 46180 234678 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 170214 45540 170220 45552
rect 3476 45512 170220 45540
rect 3476 45500 3482 45512
rect 170214 45500 170220 45512
rect 170272 45500 170278 45552
rect 152734 44956 152740 45008
rect 152792 44996 152798 45008
rect 398926 44996 398932 45008
rect 152792 44968 398932 44996
rect 152792 44956 152798 44968
rect 398926 44956 398932 44968
rect 398984 44956 398990 45008
rect 95142 44888 95148 44940
rect 95200 44928 95206 44940
rect 129090 44928 129096 44940
rect 95200 44900 129096 44928
rect 95200 44888 95206 44900
rect 129090 44888 129096 44900
rect 129148 44888 129154 44940
rect 156874 44888 156880 44940
rect 156932 44928 156938 44940
rect 447410 44928 447416 44940
rect 156932 44900 447416 44928
rect 156932 44888 156938 44900
rect 447410 44888 447416 44900
rect 447468 44888 447474 44940
rect 64322 44820 64328 44872
rect 64380 44860 64386 44872
rect 126514 44860 126520 44872
rect 64380 44832 126520 44860
rect 64380 44820 64386 44832
rect 126514 44820 126520 44832
rect 126572 44820 126578 44872
rect 160830 44820 160836 44872
rect 160888 44860 160894 44872
rect 500586 44860 500592 44872
rect 160888 44832 500592 44860
rect 160888 44820 160894 44832
rect 500586 44820 500592 44832
rect 500644 44820 500650 44872
rect 137462 43596 137468 43648
rect 137520 43636 137526 43648
rect 197906 43636 197912 43648
rect 137520 43608 197912 43636
rect 137520 43596 137526 43608
rect 197906 43596 197912 43608
rect 197964 43596 197970 43648
rect 155310 43528 155316 43580
rect 155368 43568 155374 43580
rect 434438 43568 434444 43580
rect 155368 43540 434444 43568
rect 155368 43528 155374 43540
rect 434438 43528 434444 43540
rect 434496 43528 434502 43580
rect 159542 43460 159548 43512
rect 159600 43500 159606 43512
rect 481726 43500 481732 43512
rect 159600 43472 481732 43500
rect 159600 43460 159606 43472
rect 481726 43460 481732 43472
rect 481784 43460 481790 43512
rect 133414 43392 133420 43444
rect 133472 43432 133478 43444
rect 144730 43432 144736 43444
rect 133472 43404 144736 43432
rect 133472 43392 133478 43404
rect 144730 43392 144736 43404
rect 144788 43392 144794 43444
rect 162210 43392 162216 43444
rect 162268 43432 162274 43444
rect 514754 43432 514760 43444
rect 162268 43404 514760 43432
rect 162268 43392 162274 43404
rect 514754 43392 514760 43404
rect 514812 43392 514818 43444
rect 132126 42712 132132 42764
rect 132184 42752 132190 42764
rect 132954 42752 132960 42764
rect 132184 42724 132960 42752
rect 132184 42712 132190 42724
rect 132954 42712 132960 42724
rect 133012 42712 133018 42764
rect 138842 42236 138848 42288
rect 138900 42276 138906 42288
rect 212166 42276 212172 42288
rect 138900 42248 212172 42276
rect 138900 42236 138906 42248
rect 212166 42236 212172 42248
rect 212224 42236 212230 42288
rect 149974 42168 149980 42220
rect 150032 42208 150038 42220
rect 361114 42208 361120 42220
rect 150032 42180 361120 42208
rect 150032 42168 150038 42180
rect 361114 42168 361120 42180
rect 361172 42168 361178 42220
rect 152826 42100 152832 42152
rect 152884 42140 152890 42152
rect 402514 42140 402520 42152
rect 152884 42112 402520 42140
rect 152884 42100 152890 42112
rect 402514 42100 402520 42112
rect 402572 42100 402578 42152
rect 162302 42032 162308 42084
rect 162360 42072 162366 42084
rect 525426 42072 525432 42084
rect 162360 42044 525432 42072
rect 162360 42032 162366 42044
rect 525426 42032 525432 42044
rect 525484 42032 525490 42084
rect 138934 40876 138940 40928
rect 138992 40916 138998 40928
rect 215662 40916 215668 40928
rect 138992 40888 215668 40916
rect 138992 40876 138998 40888
rect 215662 40876 215668 40888
rect 215720 40876 215726 40928
rect 142890 40808 142896 40860
rect 142948 40848 142954 40860
rect 270034 40848 270040 40860
rect 142948 40820 270040 40848
rect 142948 40808 142954 40820
rect 270034 40808 270040 40820
rect 270092 40808 270098 40860
rect 159634 40740 159640 40792
rect 159692 40780 159698 40792
rect 486418 40780 486424 40792
rect 159692 40752 486424 40780
rect 159692 40740 159698 40752
rect 486418 40740 486424 40752
rect 486476 40740 486482 40792
rect 82078 40672 82084 40724
rect 82136 40712 82142 40724
rect 120994 40712 121000 40724
rect 82136 40684 121000 40712
rect 82136 40672 82142 40684
rect 120994 40672 121000 40684
rect 121052 40672 121058 40724
rect 134426 40672 134432 40724
rect 134484 40712 134490 40724
rect 160738 40712 160744 40724
rect 134484 40684 160744 40712
rect 134484 40672 134490 40684
rect 160738 40672 160744 40684
rect 160796 40672 160802 40724
rect 160922 40672 160928 40724
rect 160980 40712 160986 40724
rect 499390 40712 499396 40724
rect 160980 40684 499396 40712
rect 160980 40672 160986 40684
rect 499390 40672 499396 40684
rect 499448 40672 499454 40724
rect 135806 39516 135812 39568
rect 135864 39556 135870 39568
rect 183738 39556 183744 39568
rect 135864 39528 183744 39556
rect 135864 39516 135870 39528
rect 183738 39516 183744 39528
rect 183796 39516 183802 39568
rect 143810 39448 143816 39500
rect 143868 39488 143874 39500
rect 286594 39488 286600 39500
rect 143868 39460 286600 39488
rect 143868 39448 143874 39460
rect 286594 39448 286600 39460
rect 286652 39448 286658 39500
rect 161014 39380 161020 39432
rect 161072 39420 161078 39432
rect 506474 39420 506480 39432
rect 161072 39392 506480 39420
rect 161072 39380 161078 39392
rect 506474 39380 506480 39392
rect 506532 39380 506538 39432
rect 163682 39312 163688 39364
rect 163740 39352 163746 39364
rect 543182 39352 543188 39364
rect 163740 39324 543188 39352
rect 163740 39312 163746 39324
rect 543182 39312 543188 39324
rect 543240 39312 543246 39364
rect 137554 38088 137560 38140
rect 137612 38128 137618 38140
rect 206186 38128 206192 38140
rect 137612 38100 206192 38128
rect 137612 38088 137618 38100
rect 206186 38088 206192 38100
rect 206244 38088 206250 38140
rect 145742 38020 145748 38072
rect 145800 38060 145806 38072
rect 300762 38060 300768 38072
rect 145800 38032 300768 38060
rect 145800 38020 145806 38032
rect 300762 38020 300768 38032
rect 300820 38020 300826 38072
rect 153838 37952 153844 38004
rect 153896 37992 153902 38004
rect 362310 37992 362316 38004
rect 153896 37964 362316 37992
rect 153896 37952 153902 37964
rect 362310 37952 362316 37964
rect 362368 37952 362374 38004
rect 166626 37884 166632 37936
rect 166684 37924 166690 37936
rect 573910 37924 573916 37936
rect 166684 37896 573916 37924
rect 166684 37884 166690 37896
rect 573910 37884 573916 37896
rect 573968 37884 573974 37936
rect 141418 36660 141424 36712
rect 141476 36700 141482 36712
rect 259454 36700 259460 36712
rect 141476 36672 259460 36700
rect 141476 36660 141482 36672
rect 259454 36660 259460 36672
rect 259512 36660 259518 36712
rect 134794 36592 134800 36644
rect 134852 36632 134858 36644
rect 156690 36632 156696 36644
rect 134852 36604 156696 36632
rect 134852 36592 134858 36604
rect 156690 36592 156696 36604
rect 156748 36592 156754 36644
rect 168282 36592 168288 36644
rect 168340 36632 168346 36644
rect 429654 36632 429660 36644
rect 168340 36604 429660 36632
rect 168340 36592 168346 36604
rect 429654 36592 429660 36604
rect 429712 36592 429718 36644
rect 155402 36524 155408 36576
rect 155460 36564 155466 36576
rect 432046 36564 432052 36576
rect 155460 36536 432052 36564
rect 155460 36524 155466 36536
rect 432046 36524 432052 36536
rect 432104 36524 432110 36576
rect 142982 35368 142988 35420
rect 143040 35408 143046 35420
rect 272426 35408 272432 35420
rect 143040 35380 272432 35408
rect 143040 35368 143046 35380
rect 272426 35368 272432 35380
rect 272484 35368 272490 35420
rect 147030 35300 147036 35352
rect 147088 35340 147094 35352
rect 319714 35340 319720 35352
rect 147088 35312 319720 35340
rect 147088 35300 147094 35312
rect 319714 35300 319720 35312
rect 319772 35300 319778 35352
rect 169202 35232 169208 35284
rect 169260 35272 169266 35284
rect 465166 35272 465172 35284
rect 169260 35244 465172 35272
rect 169260 35232 169266 35244
rect 465166 35232 465172 35244
rect 465224 35232 465230 35284
rect 161106 35164 161112 35216
rect 161164 35204 161170 35216
rect 495894 35204 495900 35216
rect 161164 35176 495900 35204
rect 161164 35164 161170 35176
rect 495894 35164 495900 35176
rect 495952 35164 495958 35216
rect 143074 33872 143080 33924
rect 143132 33912 143138 33924
rect 273622 33912 273628 33924
rect 143132 33884 273628 33912
rect 143132 33872 143138 33884
rect 273622 33872 273628 33884
rect 273680 33872 273686 33924
rect 155494 33804 155500 33856
rect 155552 33844 155558 33856
rect 424962 33844 424968 33856
rect 155552 33816 424968 33844
rect 155552 33804 155558 33816
rect 424962 33804 424968 33816
rect 425020 33804 425026 33856
rect 162394 33736 162400 33788
rect 162452 33776 162458 33788
rect 517146 33776 517152 33788
rect 162452 33748 517152 33776
rect 162452 33736 162458 33748
rect 517146 33736 517152 33748
rect 517204 33736 517210 33788
rect 139026 32648 139032 32700
rect 139084 32688 139090 32700
rect 219250 32688 219256 32700
rect 139084 32660 219256 32688
rect 139084 32648 139090 32660
rect 219250 32648 219256 32660
rect 219308 32648 219314 32700
rect 144270 32580 144276 32632
rect 144328 32620 144334 32632
rect 293678 32620 293684 32632
rect 144328 32592 293684 32620
rect 144328 32580 144334 32592
rect 293678 32580 293684 32592
rect 293736 32580 293742 32632
rect 148594 32512 148600 32564
rect 148652 32552 148658 32564
rect 337470 32552 337476 32564
rect 148652 32524 337476 32552
rect 148652 32512 148658 32524
rect 337470 32512 337476 32524
rect 337528 32512 337534 32564
rect 162578 32444 162584 32496
rect 162636 32484 162642 32496
rect 518342 32484 518348 32496
rect 162636 32456 518348 32484
rect 162636 32444 162642 32456
rect 518342 32444 518348 32456
rect 518400 32444 518406 32496
rect 133506 32376 133512 32428
rect 133564 32416 133570 32428
rect 142430 32416 142436 32428
rect 133564 32388 142436 32416
rect 133564 32376 133570 32388
rect 142430 32376 142436 32388
rect 142488 32376 142494 32428
rect 162486 32376 162492 32428
rect 162544 32416 162550 32428
rect 520734 32416 520740 32428
rect 162544 32388 520740 32416
rect 162544 32376 162550 32388
rect 520734 32376 520740 32388
rect 520792 32376 520798 32428
rect 140314 31288 140320 31340
rect 140372 31328 140378 31340
rect 233418 31328 233424 31340
rect 140372 31300 233424 31328
rect 140372 31288 140378 31300
rect 233418 31288 233424 31300
rect 233476 31288 233482 31340
rect 150066 31220 150072 31272
rect 150124 31260 150130 31272
rect 357526 31260 357532 31272
rect 150124 31232 357532 31260
rect 150124 31220 150130 31232
rect 357526 31220 357532 31232
rect 357584 31220 357590 31272
rect 159726 31152 159732 31204
rect 159784 31192 159790 31204
rect 485222 31192 485228 31204
rect 159784 31164 485228 31192
rect 159784 31152 159790 31164
rect 485222 31152 485228 31164
rect 485280 31152 485286 31204
rect 163774 31084 163780 31136
rect 163832 31124 163838 31136
rect 536098 31124 536104 31136
rect 163832 31096 536104 31124
rect 163832 31084 163838 31096
rect 536098 31084 536104 31096
rect 536156 31084 536162 31136
rect 134886 31016 134892 31068
rect 134944 31056 134950 31068
rect 162118 31056 162124 31068
rect 134944 31028 162124 31056
rect 134944 31016 134950 31028
rect 162118 31016 162124 31028
rect 162176 31016 162182 31068
rect 165246 31016 165252 31068
rect 165304 31056 165310 31068
rect 549070 31056 549076 31068
rect 165304 31028 549076 31056
rect 165304 31016 165310 31028
rect 549070 31016 549076 31028
rect 549128 31016 549134 31068
rect 134978 29724 134984 29776
rect 135036 29764 135042 29776
rect 158070 29764 158076 29776
rect 135036 29736 158076 29764
rect 135036 29724 135042 29736
rect 158070 29724 158076 29736
rect 158128 29724 158134 29776
rect 156966 29656 156972 29708
rect 157024 29696 157030 29708
rect 454494 29696 454500 29708
rect 157024 29668 454500 29696
rect 157024 29656 157030 29668
rect 454494 29656 454500 29668
rect 454552 29656 454558 29708
rect 157334 29588 157340 29640
rect 157392 29628 157398 29640
rect 460382 29628 460388 29640
rect 157392 29600 460388 29628
rect 157392 29588 157398 29600
rect 460382 29588 460388 29600
rect 460440 29588 460446 29640
rect 139118 28568 139124 28620
rect 139176 28608 139182 28620
rect 223942 28608 223948 28620
rect 139176 28580 223948 28608
rect 139176 28568 139182 28580
rect 223942 28568 223948 28580
rect 224000 28568 224006 28620
rect 143166 28500 143172 28552
rect 143224 28540 143230 28552
rect 268838 28540 268844 28552
rect 143224 28512 268844 28540
rect 143224 28500 143230 28512
rect 268838 28500 268844 28512
rect 268896 28500 268902 28552
rect 151262 28432 151268 28484
rect 151320 28472 151326 28484
rect 372890 28472 372896 28484
rect 151320 28444 372896 28472
rect 151320 28432 151326 28444
rect 372890 28432 372896 28444
rect 372948 28432 372954 28484
rect 155954 28364 155960 28416
rect 156012 28404 156018 28416
rect 449802 28404 449808 28416
rect 156012 28376 449808 28404
rect 156012 28364 156018 28376
rect 449802 28364 449808 28376
rect 449860 28364 449866 28416
rect 159818 28296 159824 28348
rect 159876 28336 159882 28348
rect 488810 28336 488816 28348
rect 159876 28308 488816 28336
rect 159876 28296 159882 28308
rect 488810 28296 488816 28308
rect 488868 28296 488874 28348
rect 166718 28228 166724 28280
rect 166776 28268 166782 28280
rect 566826 28268 566832 28280
rect 166776 28240 566832 28268
rect 166776 28228 166782 28240
rect 566826 28228 566832 28240
rect 566884 28228 566890 28280
rect 149698 27072 149704 27124
rect 149756 27112 149762 27124
rect 315022 27112 315028 27124
rect 149756 27084 315028 27112
rect 149756 27072 149762 27084
rect 315022 27072 315028 27084
rect 315080 27072 315086 27124
rect 151354 27004 151360 27056
rect 151412 27044 151418 27056
rect 379974 27044 379980 27056
rect 151412 27016 379980 27044
rect 151412 27004 151418 27016
rect 379974 27004 379980 27016
rect 380032 27004 380038 27056
rect 160370 26936 160376 26988
rect 160428 26976 160434 26988
rect 507670 26976 507676 26988
rect 160428 26948 507676 26976
rect 160428 26936 160434 26948
rect 507670 26936 507676 26948
rect 507728 26936 507734 26988
rect 165890 26868 165896 26920
rect 165948 26908 165954 26920
rect 570322 26908 570328 26920
rect 165948 26880 570328 26908
rect 165948 26868 165954 26880
rect 570322 26868 570328 26880
rect 570380 26868 570386 26920
rect 145834 25712 145840 25764
rect 145892 25752 145898 25764
rect 304350 25752 304356 25764
rect 145892 25724 304356 25752
rect 145892 25712 145898 25724
rect 304350 25712 304356 25724
rect 304408 25712 304414 25764
rect 151446 25644 151452 25696
rect 151504 25684 151510 25696
rect 371694 25684 371700 25696
rect 151504 25656 371700 25684
rect 151504 25644 151510 25656
rect 371694 25644 371700 25656
rect 371752 25644 371758 25696
rect 160462 25576 160468 25628
rect 160520 25616 160526 25628
rect 502978 25616 502984 25628
rect 160520 25588 502984 25616
rect 160520 25576 160526 25588
rect 502978 25576 502984 25588
rect 503036 25576 503042 25628
rect 20622 25508 20628 25560
rect 20680 25548 20686 25560
rect 107010 25548 107016 25560
rect 20680 25520 107016 25548
rect 20680 25508 20686 25520
rect 107010 25508 107016 25520
rect 107068 25508 107074 25560
rect 161750 25508 161756 25560
rect 161808 25548 161814 25560
rect 521838 25548 521844 25560
rect 161808 25520 521844 25548
rect 161808 25508 161814 25520
rect 521838 25508 521844 25520
rect 521896 25508 521902 25560
rect 140406 24420 140412 24472
rect 140464 24460 140470 24472
rect 237006 24460 237012 24472
rect 140464 24432 237012 24460
rect 140464 24420 140470 24432
rect 237006 24420 237012 24432
rect 237064 24420 237070 24472
rect 147122 24352 147128 24404
rect 147180 24392 147186 24404
rect 318518 24392 318524 24404
rect 147180 24364 318524 24392
rect 147180 24352 147186 24364
rect 318518 24352 318524 24364
rect 318576 24352 318582 24404
rect 152918 24284 152924 24336
rect 152976 24324 152982 24336
rect 389450 24324 389456 24336
rect 152976 24296 389456 24324
rect 152976 24284 152982 24296
rect 389450 24284 389456 24296
rect 389508 24284 389514 24336
rect 168190 24216 168196 24268
rect 168248 24256 168254 24268
rect 408402 24256 408408 24268
rect 168248 24228 408408 24256
rect 168248 24216 168254 24228
rect 408402 24216 408408 24228
rect 408460 24216 408466 24268
rect 160646 24148 160652 24200
rect 160704 24188 160710 24200
rect 510062 24188 510068 24200
rect 160704 24160 510068 24188
rect 160704 24148 160710 24160
rect 510062 24148 510068 24160
rect 510120 24148 510126 24200
rect 163866 24080 163872 24132
rect 163924 24120 163930 24132
rect 532510 24120 532516 24132
rect 163924 24092 532516 24120
rect 163924 24080 163930 24092
rect 532510 24080 532516 24092
rect 532568 24080 532574 24132
rect 144362 22856 144368 22908
rect 144420 22896 144426 22908
rect 287790 22896 287796 22908
rect 144420 22868 287796 22896
rect 144420 22856 144426 22868
rect 287790 22856 287796 22868
rect 287848 22856 287854 22908
rect 168098 22788 168104 22840
rect 168156 22828 168162 22840
rect 401318 22828 401324 22840
rect 168156 22800 401324 22828
rect 168156 22788 168162 22800
rect 401318 22788 401324 22800
rect 401376 22788 401382 22840
rect 161474 22720 161480 22772
rect 161532 22760 161538 22772
rect 513558 22760 513564 22772
rect 161532 22732 513564 22760
rect 161532 22720 161538 22732
rect 513558 22720 513564 22732
rect 513616 22720 513622 22772
rect 140498 21632 140504 21684
rect 140556 21672 140562 21684
rect 231026 21672 231032 21684
rect 140556 21644 231032 21672
rect 140556 21632 140562 21644
rect 231026 21632 231032 21644
rect 231084 21632 231090 21684
rect 148778 21564 148784 21616
rect 148836 21604 148842 21616
rect 340966 21604 340972 21616
rect 148836 21576 340972 21604
rect 148836 21564 148842 21576
rect 340966 21564 340972 21576
rect 341024 21564 341030 21616
rect 148686 21496 148692 21548
rect 148744 21536 148750 21548
rect 344554 21536 344560 21548
rect 148744 21508 344560 21536
rect 148744 21496 148750 21508
rect 344554 21496 344560 21508
rect 344612 21496 344618 21548
rect 149146 21428 149152 21480
rect 149204 21468 149210 21480
rect 358722 21468 358728 21480
rect 149204 21440 358728 21468
rect 149204 21428 149210 21440
rect 358722 21428 358728 21440
rect 358780 21428 358786 21480
rect 133598 21360 133604 21412
rect 133656 21400 133662 21412
rect 148318 21400 148324 21412
rect 133656 21372 148324 21400
rect 133656 21360 133662 21372
rect 148318 21360 148324 21372
rect 148376 21360 148382 21412
rect 149238 21360 149244 21412
rect 149296 21400 149302 21412
rect 365806 21400 365812 21412
rect 149296 21372 365812 21400
rect 149296 21360 149302 21372
rect 365806 21360 365812 21372
rect 365864 21360 365870 21412
rect 143258 20204 143264 20256
rect 143316 20244 143322 20256
rect 266538 20244 266544 20256
rect 143316 20216 266544 20244
rect 143316 20204 143322 20216
rect 266538 20204 266544 20216
rect 266596 20204 266602 20256
rect 144546 20136 144552 20188
rect 144604 20176 144610 20188
rect 284294 20176 284300 20188
rect 144604 20148 284300 20176
rect 144604 20136 144610 20148
rect 284294 20136 284300 20148
rect 284352 20136 284358 20188
rect 144454 20068 144460 20120
rect 144512 20108 144518 20120
rect 294874 20108 294880 20120
rect 144512 20080 294880 20108
rect 144512 20068 144518 20080
rect 294874 20068 294880 20080
rect 294932 20068 294938 20120
rect 159358 20000 159364 20052
rect 159416 20040 159422 20052
rect 383562 20040 383568 20052
rect 159416 20012 383568 20040
rect 159416 20000 159422 20012
rect 383562 20000 383568 20012
rect 383620 20000 383626 20052
rect 169110 19932 169116 19984
rect 169168 19972 169174 19984
rect 450906 19972 450912 19984
rect 169168 19944 450912 19972
rect 169168 19932 169174 19944
rect 450906 19932 450912 19944
rect 450964 19932 450970 19984
rect 137646 18776 137652 18828
rect 137704 18816 137710 18828
rect 202690 18816 202696 18828
rect 137704 18788 202696 18816
rect 137704 18776 137710 18788
rect 202690 18776 202696 18788
rect 202748 18776 202754 18828
rect 139670 18708 139676 18760
rect 139728 18748 139734 18760
rect 238110 18748 238116 18760
rect 139728 18720 238116 18748
rect 139728 18708 139734 18720
rect 238110 18708 238116 18720
rect 238168 18708 238174 18760
rect 151538 18640 151544 18692
rect 151596 18680 151602 18692
rect 376478 18680 376484 18692
rect 151596 18652 376484 18680
rect 151596 18640 151602 18652
rect 376478 18640 376484 18652
rect 376536 18640 376542 18692
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 116854 18612 116860 18624
rect 11204 18584 116860 18612
rect 11204 18572 11210 18584
rect 116854 18572 116860 18584
rect 116912 18572 116918 18624
rect 166074 18572 166080 18624
rect 166132 18612 166138 18624
rect 571518 18612 571524 18624
rect 166132 18584 571524 18612
rect 166132 18572 166138 18584
rect 571518 18572 571524 18584
rect 571576 18572 571582 18624
rect 138290 17484 138296 17536
rect 138348 17524 138354 17536
rect 220446 17524 220452 17536
rect 138348 17496 220452 17524
rect 138348 17484 138354 17496
rect 220446 17484 220452 17496
rect 220504 17484 220510 17536
rect 168006 17416 168012 17468
rect 168064 17456 168070 17468
rect 443822 17456 443828 17468
rect 168064 17428 443828 17456
rect 168064 17416 168070 17428
rect 443822 17416 443828 17428
rect 443880 17416 443886 17468
rect 157610 17348 157616 17400
rect 157668 17388 157674 17400
rect 463970 17388 463976 17400
rect 157668 17360 463976 17388
rect 157668 17348 157674 17360
rect 463970 17348 463976 17360
rect 464028 17348 464034 17400
rect 157426 17280 157432 17332
rect 157484 17320 157490 17332
rect 467466 17320 467472 17332
rect 157484 17292 467472 17320
rect 157484 17280 157490 17292
rect 467466 17280 467472 17292
rect 467524 17280 467530 17332
rect 43070 17212 43076 17264
rect 43128 17252 43134 17264
rect 109678 17252 109684 17264
rect 43128 17224 109684 17252
rect 43128 17212 43134 17224
rect 109678 17212 109684 17224
rect 109736 17212 109742 17264
rect 132586 17212 132592 17264
rect 132644 17252 132650 17264
rect 151078 17252 151084 17264
rect 132644 17224 151084 17252
rect 132644 17212 132650 17224
rect 151078 17212 151084 17224
rect 151136 17212 151142 17264
rect 157794 17212 157800 17264
rect 157852 17252 157858 17264
rect 471054 17252 471060 17264
rect 157852 17224 471060 17252
rect 157852 17212 157858 17224
rect 471054 17212 471060 17224
rect 471112 17212 471118 17264
rect 138474 16124 138480 16176
rect 138532 16164 138538 16176
rect 222746 16164 222752 16176
rect 138532 16136 222752 16164
rect 138532 16124 138538 16136
rect 222746 16124 222752 16136
rect 222804 16124 222810 16176
rect 147214 16056 147220 16108
rect 147272 16096 147278 16108
rect 323302 16096 323308 16108
rect 147272 16068 323308 16096
rect 147272 16056 147278 16068
rect 323302 16056 323308 16068
rect 323360 16056 323366 16108
rect 150710 15988 150716 16040
rect 150768 16028 150774 16040
rect 375282 16028 375288 16040
rect 150768 16000 375288 16028
rect 150768 15988 150774 16000
rect 375282 15988 375288 16000
rect 375340 15988 375346 16040
rect 150526 15920 150532 15972
rect 150584 15960 150590 15972
rect 378870 15960 378876 15972
rect 150584 15932 378876 15960
rect 150584 15920 150590 15932
rect 378870 15920 378876 15932
rect 378928 15920 378934 15972
rect 35986 15852 35992 15904
rect 36044 15892 36050 15904
rect 113910 15892 113916 15904
rect 36044 15864 113916 15892
rect 36044 15852 36050 15864
rect 113910 15852 113916 15864
rect 113968 15852 113974 15904
rect 152182 15852 152188 15904
rect 152240 15892 152246 15904
rect 393038 15892 393044 15904
rect 152240 15864 393044 15892
rect 152240 15852 152246 15864
rect 393038 15852 393044 15864
rect 393096 15852 393102 15904
rect 143350 14696 143356 14748
rect 143408 14736 143414 14748
rect 276014 14736 276020 14748
rect 143408 14708 276020 14736
rect 143408 14696 143414 14708
rect 276014 14696 276020 14708
rect 276072 14696 276078 14748
rect 144638 14628 144644 14680
rect 144696 14668 144702 14680
rect 290182 14668 290188 14680
rect 144696 14640 290188 14668
rect 144696 14628 144702 14640
rect 290182 14628 290188 14640
rect 290240 14628 290246 14680
rect 148134 14560 148140 14612
rect 148192 14600 148198 14612
rect 336274 14600 336280 14612
rect 148192 14572 336280 14600
rect 148192 14560 148198 14572
rect 336274 14560 336280 14572
rect 336332 14560 336338 14612
rect 167914 14492 167920 14544
rect 167972 14532 167978 14544
rect 422570 14532 422576 14544
rect 167972 14504 422576 14532
rect 167972 14492 167978 14504
rect 422570 14492 422576 14504
rect 422628 14492 422634 14544
rect 28902 14424 28908 14476
rect 28960 14464 28966 14476
rect 118142 14464 118148 14476
rect 28960 14436 118148 14464
rect 28960 14424 28966 14436
rect 118142 14424 118148 14436
rect 118200 14424 118206 14476
rect 154206 14424 154212 14476
rect 154264 14464 154270 14476
rect 414290 14464 414296 14476
rect 154264 14436 414296 14464
rect 154264 14424 154270 14436
rect 414290 14424 414296 14436
rect 414348 14424 414354 14476
rect 139854 13336 139860 13388
rect 139912 13376 139918 13388
rect 240502 13376 240508 13388
rect 139912 13348 240508 13376
rect 139912 13336 139918 13348
rect 240502 13336 240508 13348
rect 240560 13336 240566 13388
rect 147306 13268 147312 13320
rect 147364 13308 147370 13320
rect 325602 13308 325608 13320
rect 147364 13280 325608 13308
rect 147364 13268 147370 13280
rect 325602 13268 325608 13280
rect 325660 13268 325666 13320
rect 154298 13200 154304 13252
rect 154356 13240 154362 13252
rect 410794 13240 410800 13252
rect 154356 13212 410800 13240
rect 154356 13200 154362 13212
rect 410794 13200 410800 13212
rect 410852 13200 410858 13252
rect 155586 13132 155592 13184
rect 155644 13172 155650 13184
rect 426158 13172 426164 13184
rect 155644 13144 426164 13172
rect 155644 13132 155650 13144
rect 426158 13132 426164 13144
rect 426216 13132 426222 13184
rect 85666 13064 85672 13116
rect 85724 13104 85730 13116
rect 120902 13104 120908 13116
rect 85724 13076 120908 13104
rect 85724 13064 85730 13076
rect 120902 13064 120908 13076
rect 120960 13064 120966 13116
rect 133966 13064 133972 13116
rect 134024 13104 134030 13116
rect 153838 13104 153844 13116
rect 134024 13076 153844 13104
rect 134024 13064 134030 13076
rect 153838 13064 153844 13076
rect 153896 13064 153902 13116
rect 165338 13064 165344 13116
rect 165396 13104 165402 13116
rect 550266 13104 550272 13116
rect 165396 13076 550272 13104
rect 165396 13064 165402 13076
rect 550266 13064 550272 13076
rect 550324 13064 550330 13116
rect 132218 12384 132224 12436
rect 132276 12424 132282 12436
rect 133138 12424 133144 12436
rect 132276 12396 133144 12424
rect 132276 12384 132282 12396
rect 133138 12384 133144 12396
rect 133196 12384 133202 12436
rect 167822 11772 167828 11824
rect 167880 11812 167886 11824
rect 415486 11812 415492 11824
rect 167880 11784 415492 11812
rect 167880 11772 167886 11784
rect 415486 11772 415492 11784
rect 415544 11772 415550 11824
rect 158990 11704 158996 11756
rect 159048 11744 159054 11756
rect 482830 11744 482836 11756
rect 159048 11716 482836 11744
rect 159048 11704 159054 11716
rect 482830 11704 482836 11716
rect 482888 11704 482894 11756
rect 147398 10480 147404 10532
rect 147456 10520 147462 10532
rect 329190 10520 329196 10532
rect 147456 10492 329196 10520
rect 147456 10480 147462 10492
rect 329190 10480 329196 10492
rect 329248 10480 329254 10532
rect 155678 10412 155684 10464
rect 155736 10452 155742 10464
rect 435542 10452 435548 10464
rect 155736 10424 435548 10452
rect 155736 10412 155742 10424
rect 435542 10412 435548 10424
rect 435600 10412 435606 10464
rect 46658 10344 46664 10396
rect 46716 10384 46722 10396
rect 125502 10384 125508 10396
rect 46716 10356 125508 10384
rect 46716 10344 46722 10356
rect 125502 10344 125508 10356
rect 125560 10344 125566 10396
rect 169018 10344 169024 10396
rect 169076 10384 169082 10396
rect 458082 10384 458088 10396
rect 169076 10356 458088 10384
rect 169076 10344 169082 10356
rect 458082 10344 458088 10356
rect 458140 10344 458146 10396
rect 19426 10276 19432 10328
rect 19484 10316 19490 10328
rect 118050 10316 118056 10328
rect 19484 10288 118056 10316
rect 19484 10276 19490 10288
rect 118050 10276 118056 10288
rect 118108 10276 118114 10328
rect 163958 10276 163964 10328
rect 164016 10316 164022 10328
rect 534902 10316 534908 10328
rect 164016 10288 534908 10316
rect 164016 10276 164022 10288
rect 534902 10276 534908 10288
rect 534960 10276 534966 10328
rect 145926 9256 145932 9308
rect 145984 9296 145990 9308
rect 309042 9296 309048 9308
rect 145984 9268 309048 9296
rect 145984 9256 145990 9268
rect 309042 9256 309048 9268
rect 309100 9256 309106 9308
rect 145098 9188 145104 9240
rect 145156 9228 145162 9240
rect 312630 9228 312636 9240
rect 145156 9200 312636 9228
rect 145156 9188 145162 9200
rect 312630 9188 312636 9200
rect 312688 9188 312694 9240
rect 149422 9120 149428 9172
rect 149480 9160 149486 9172
rect 364610 9160 364616 9172
rect 149480 9132 364616 9160
rect 149480 9120 149486 9132
rect 364610 9120 364616 9132
rect 364668 9120 364674 9172
rect 154390 9052 154396 9104
rect 154448 9092 154454 9104
rect 411898 9092 411904 9104
rect 154448 9064 411904 9092
rect 154448 9052 154454 9064
rect 411898 9052 411904 9064
rect 411956 9052 411962 9104
rect 159174 8984 159180 9036
rect 159232 9024 159238 9036
rect 478138 9024 478144 9036
rect 159232 8996 478144 9024
rect 159232 8984 159238 8996
rect 478138 8984 478144 8996
rect 478196 8984 478202 9036
rect 96246 8916 96252 8968
rect 96304 8956 96310 8968
rect 128906 8956 128912 8968
rect 96304 8928 128912 8956
rect 96304 8916 96310 8928
rect 128906 8916 128912 8928
rect 128964 8916 128970 8968
rect 164050 8916 164056 8968
rect 164108 8956 164114 8968
rect 531314 8956 531320 8968
rect 164108 8928 531320 8956
rect 164108 8916 164114 8928
rect 531314 8916 531320 8928
rect 531372 8916 531378 8968
rect 471238 8236 471244 8288
rect 471296 8276 471302 8288
rect 479334 8276 479340 8288
rect 471296 8248 479340 8276
rect 471296 8236 471302 8248
rect 479334 8236 479340 8248
rect 479392 8236 479398 8288
rect 142154 7760 142160 7812
rect 142212 7800 142218 7812
rect 265342 7800 265348 7812
rect 142212 7772 265348 7800
rect 142212 7760 142218 7772
rect 265342 7760 265348 7772
rect 265400 7760 265406 7812
rect 147950 7692 147956 7744
rect 148008 7732 148014 7744
rect 339862 7732 339868 7744
rect 148008 7704 339868 7732
rect 148008 7692 148014 7704
rect 339862 7692 339868 7704
rect 339920 7692 339926 7744
rect 50154 7624 50160 7676
rect 50212 7664 50218 7676
rect 125410 7664 125416 7676
rect 50212 7636 125416 7664
rect 50212 7624 50218 7636
rect 125410 7624 125416 7636
rect 125468 7624 125474 7676
rect 155770 7624 155776 7676
rect 155828 7664 155834 7676
rect 428458 7664 428464 7676
rect 155828 7636 428464 7664
rect 155828 7624 155834 7636
rect 428458 7624 428464 7636
rect 428516 7624 428522 7676
rect 24210 7556 24216 7608
rect 24268 7596 24274 7608
rect 116762 7596 116768 7608
rect 24268 7568 116768 7596
rect 24268 7556 24274 7568
rect 116762 7556 116768 7568
rect 116820 7556 116826 7608
rect 163222 7556 163228 7608
rect 163280 7596 163286 7608
rect 541986 7596 541992 7608
rect 163280 7568 541992 7596
rect 163280 7556 163286 7568
rect 541986 7556 541992 7568
rect 542044 7556 542050 7608
rect 141786 6808 141792 6860
rect 141844 6848 141850 6860
rect 248782 6848 248788 6860
rect 141844 6820 248788 6848
rect 141844 6808 141850 6820
rect 248782 6808 248788 6820
rect 248840 6808 248846 6860
rect 141510 6740 141516 6792
rect 141568 6780 141574 6792
rect 252370 6780 252376 6792
rect 141568 6752 252376 6780
rect 141568 6740 141574 6752
rect 252370 6740 252376 6752
rect 252428 6740 252434 6792
rect 141602 6672 141608 6724
rect 141660 6712 141666 6724
rect 254670 6712 254676 6724
rect 141660 6684 254676 6712
rect 141660 6672 141666 6684
rect 254670 6672 254676 6684
rect 254728 6672 254734 6724
rect 141878 6604 141884 6656
rect 141936 6644 141942 6656
rect 258258 6644 258264 6656
rect 141936 6616 258264 6644
rect 141936 6604 141942 6616
rect 258258 6604 258264 6616
rect 258316 6604 258322 6656
rect 141694 6536 141700 6588
rect 141752 6576 141758 6588
rect 261754 6576 261760 6588
rect 141752 6548 261760 6576
rect 141752 6536 141758 6548
rect 261754 6536 261760 6548
rect 261812 6536 261818 6588
rect 2774 6468 2780 6520
rect 2832 6508 2838 6520
rect 4798 6508 4804 6520
rect 2832 6480 4804 6508
rect 2832 6468 2838 6480
rect 4798 6468 4804 6480
rect 4856 6468 4862 6520
rect 145006 6468 145012 6520
rect 145064 6508 145070 6520
rect 301958 6508 301964 6520
rect 145064 6480 301964 6508
rect 145064 6468 145070 6480
rect 301958 6468 301964 6480
rect 302016 6468 302022 6520
rect 145374 6400 145380 6452
rect 145432 6440 145438 6452
rect 305546 6440 305552 6452
rect 145432 6412 305552 6440
rect 145432 6400 145438 6412
rect 305546 6400 305552 6412
rect 305604 6400 305610 6452
rect 153194 6332 153200 6384
rect 153252 6372 153258 6384
rect 417878 6372 417884 6384
rect 153252 6344 417884 6372
rect 153252 6332 153258 6344
rect 417878 6332 417884 6344
rect 417936 6332 417942 6384
rect 154666 6264 154672 6316
rect 154724 6304 154730 6316
rect 433242 6304 433248 6316
rect 154724 6276 433248 6304
rect 154724 6264 154730 6276
rect 433242 6264 433248 6276
rect 433300 6264 433306 6316
rect 78582 6196 78588 6248
rect 78640 6236 78646 6248
rect 127434 6236 127440 6248
rect 78640 6208 127440 6236
rect 78640 6196 78646 6208
rect 127434 6196 127440 6208
rect 127492 6196 127498 6248
rect 132402 6196 132408 6248
rect 132460 6236 132466 6248
rect 137646 6236 137652 6248
rect 132460 6208 137652 6236
rect 132460 6196 132466 6208
rect 137646 6196 137652 6208
rect 137704 6196 137710 6248
rect 164602 6196 164608 6248
rect 164660 6236 164666 6248
rect 556154 6236 556160 6248
rect 164660 6208 556160 6236
rect 164660 6196 164666 6208
rect 556154 6196 556160 6208
rect 556212 6196 556218 6248
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 122190 6168 122196 6180
rect 6512 6140 122196 6168
rect 6512 6128 6518 6140
rect 122190 6128 122196 6140
rect 122248 6128 122254 6180
rect 122282 6128 122288 6180
rect 122340 6168 122346 6180
rect 127618 6168 127624 6180
rect 122340 6140 127624 6168
rect 122340 6128 122346 6140
rect 127618 6128 127624 6140
rect 127676 6128 127682 6180
rect 132770 6128 132776 6180
rect 132828 6168 132834 6180
rect 151814 6168 151820 6180
rect 132828 6140 151820 6168
rect 132828 6128 132834 6140
rect 151814 6128 151820 6140
rect 151872 6128 151878 6180
rect 164786 6128 164792 6180
rect 164844 6168 164850 6180
rect 557350 6168 557356 6180
rect 164844 6140 557356 6168
rect 164844 6128 164850 6140
rect 557350 6128 557356 6140
rect 557408 6128 557414 6180
rect 136818 6060 136824 6112
rect 136876 6100 136882 6112
rect 205082 6100 205088 6112
rect 136876 6072 205088 6100
rect 136876 6060 136882 6072
rect 205082 6060 205088 6072
rect 205140 6060 205146 6112
rect 137738 5992 137744 6044
rect 137796 6032 137802 6044
rect 195606 6032 195612 6044
rect 137796 6004 195612 6032
rect 137796 5992 137802 6004
rect 195606 5992 195612 6004
rect 195664 5992 195670 6044
rect 132310 5516 132316 5568
rect 132368 5556 132374 5568
rect 133782 5556 133788 5568
rect 132368 5528 133788 5556
rect 132368 5516 132374 5528
rect 133782 5516 133788 5528
rect 133840 5516 133846 5568
rect 137002 5108 137008 5160
rect 137060 5148 137066 5160
rect 199102 5148 199108 5160
rect 137060 5120 199108 5148
rect 137060 5108 137066 5120
rect 199102 5108 199108 5120
rect 199160 5108 199166 5160
rect 146478 5040 146484 5092
rect 146536 5080 146542 5092
rect 322106 5080 322112 5092
rect 146536 5052 322112 5080
rect 146536 5040 146542 5052
rect 322106 5040 322112 5052
rect 322164 5040 322170 5092
rect 147490 4972 147496 5024
rect 147548 5012 147554 5024
rect 330386 5012 330392 5024
rect 147548 4984 330392 5012
rect 147548 4972 147554 4984
rect 330386 4972 330392 4984
rect 330444 4972 330450 5024
rect 157978 4904 157984 4956
rect 158036 4944 158042 4956
rect 390646 4944 390652 4956
rect 158036 4916 390652 4944
rect 158036 4904 158042 4916
rect 390646 4904 390652 4916
rect 390704 4904 390710 4956
rect 71498 4836 71504 4888
rect 71556 4876 71562 4888
rect 120718 4876 120724 4888
rect 71556 4848 120724 4876
rect 71556 4836 71562 4848
rect 120718 4836 120724 4848
rect 120776 4836 120782 4888
rect 152366 4836 152372 4888
rect 152424 4876 152430 4888
rect 400122 4876 400128 4888
rect 152424 4848 400128 4876
rect 152424 4836 152430 4848
rect 400122 4836 400128 4848
rect 400180 4836 400186 4888
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 25498 4808 25504 4820
rect 5316 4780 25504 4808
rect 5316 4768 5322 4780
rect 25498 4768 25504 4780
rect 25556 4768 25562 4820
rect 45462 4768 45468 4820
rect 45520 4808 45526 4820
rect 125226 4808 125232 4820
rect 45520 4780 125232 4808
rect 45520 4768 45526 4780
rect 125226 4768 125232 4780
rect 125284 4768 125290 4820
rect 134518 4768 134524 4820
rect 134576 4808 134582 4820
rect 143534 4808 143540 4820
rect 134576 4780 143540 4808
rect 134576 4768 134582 4780
rect 143534 4768 143540 4780
rect 143592 4768 143598 4820
rect 166258 4768 166264 4820
rect 166316 4808 166322 4820
rect 498194 4808 498200 4820
rect 166316 4780 498200 4808
rect 166316 4768 166322 4780
rect 498194 4768 498200 4780
rect 498252 4768 498258 4820
rect 141142 4088 141148 4140
rect 141200 4128 141206 4140
rect 257062 4128 257068 4140
rect 141200 4100 257068 4128
rect 141200 4088 141206 4100
rect 257062 4088 257068 4100
rect 257120 4088 257126 4140
rect 141234 4020 141240 4072
rect 141292 4060 141298 4072
rect 260650 4060 260656 4072
rect 141292 4032 260656 4060
rect 141292 4020 141298 4032
rect 260650 4020 260656 4032
rect 260708 4020 260714 4072
rect 151078 3952 151084 4004
rect 151136 3992 151142 4004
rect 153010 3992 153016 4004
rect 151136 3964 153016 3992
rect 151136 3952 151142 3964
rect 153010 3952 153016 3964
rect 153068 3952 153074 4004
rect 160738 3952 160744 4004
rect 160796 3992 160802 4004
rect 162486 3992 162492 4004
rect 160796 3964 162492 3992
rect 160796 3952 160802 3964
rect 162486 3952 162492 3964
rect 162544 3952 162550 4004
rect 167638 3952 167644 4004
rect 167696 3992 167702 4004
rect 303154 3992 303160 4004
rect 167696 3964 303160 3992
rect 167696 3952 167702 3964
rect 303154 3952 303160 3964
rect 303212 3952 303218 4004
rect 143994 3884 144000 3936
rect 144052 3924 144058 3936
rect 292574 3924 292580 3936
rect 144052 3896 292580 3924
rect 144052 3884 144058 3896
rect 292574 3884 292580 3896
rect 292632 3884 292638 3936
rect 108114 3816 108120 3868
rect 108172 3856 108178 3868
rect 119338 3856 119344 3868
rect 108172 3828 119344 3856
rect 108172 3816 108178 3828
rect 119338 3816 119344 3828
rect 119396 3816 119402 3868
rect 170398 3816 170404 3868
rect 170456 3856 170462 3868
rect 187326 3856 187332 3868
rect 170456 3828 187332 3856
rect 170456 3816 170462 3828
rect 187326 3816 187332 3828
rect 187384 3816 187390 3868
rect 189810 3816 189816 3868
rect 189868 3856 189874 3868
rect 346946 3856 346952 3868
rect 189868 3828 346952 3856
rect 189868 3816 189874 3828
rect 346946 3816 346952 3828
rect 347004 3816 347010 3868
rect 98638 3748 98644 3800
rect 98696 3788 98702 3800
rect 111058 3788 111064 3800
rect 98696 3760 111064 3788
rect 98696 3748 98702 3760
rect 111058 3748 111064 3760
rect 111116 3748 111122 3800
rect 136174 3748 136180 3800
rect 136232 3788 136238 3800
rect 147122 3788 147128 3800
rect 136232 3760 147128 3788
rect 136232 3748 136238 3760
rect 147122 3748 147128 3760
rect 147180 3748 147186 3800
rect 156230 3748 156236 3800
rect 156288 3788 156294 3800
rect 452102 3788 452108 3800
rect 156288 3760 452108 3788
rect 156288 3748 156294 3760
rect 452102 3748 452108 3760
rect 452160 3748 452166 3800
rect 66714 3680 66720 3732
rect 66772 3720 66778 3732
rect 120810 3720 120816 3732
rect 66772 3692 120816 3720
rect 66772 3680 66778 3692
rect 120810 3680 120816 3692
rect 120868 3680 120874 3732
rect 134610 3680 134616 3732
rect 134668 3720 134674 3732
rect 145926 3720 145932 3732
rect 134668 3692 145932 3720
rect 134668 3680 134674 3692
rect 145926 3680 145932 3692
rect 145984 3680 145990 3732
rect 167730 3680 167736 3732
rect 167788 3720 167794 3732
rect 462774 3720 462780 3732
rect 167788 3692 462780 3720
rect 167788 3680 167794 3692
rect 462774 3680 462780 3692
rect 462832 3680 462838 3732
rect 51350 3612 51356 3664
rect 51408 3652 51414 3664
rect 119522 3652 119528 3664
rect 51408 3624 119528 3652
rect 51408 3612 51414 3624
rect 119522 3612 119528 3624
rect 119580 3612 119586 3664
rect 135898 3612 135904 3664
rect 135956 3652 135962 3664
rect 149514 3652 149520 3664
rect 135956 3624 149520 3652
rect 135956 3612 135962 3624
rect 149514 3612 149520 3624
rect 149572 3612 149578 3664
rect 151170 3612 151176 3664
rect 151228 3652 151234 3664
rect 155402 3652 155408 3664
rect 151228 3624 155408 3652
rect 151228 3612 151234 3624
rect 155402 3612 155408 3624
rect 155460 3612 155466 3664
rect 156414 3612 156420 3664
rect 156472 3652 156478 3664
rect 455690 3652 455696 3664
rect 156472 3624 455696 3652
rect 156472 3612 156478 3624
rect 455690 3612 455696 3624
rect 455748 3612 455754 3664
rect 475378 3612 475384 3664
rect 475436 3652 475442 3664
rect 546678 3652 546684 3664
rect 475436 3624 546684 3652
rect 475436 3612 475442 3624
rect 546678 3612 546684 3624
rect 546736 3612 546742 3664
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 119430 3584 119436 3596
rect 15988 3556 119436 3584
rect 15988 3544 15994 3556
rect 119430 3544 119436 3556
rect 119488 3544 119494 3596
rect 135990 3544 135996 3596
rect 136048 3584 136054 3596
rect 150618 3584 150624 3596
rect 136048 3556 150624 3584
rect 136048 3544 136054 3556
rect 150618 3544 150624 3556
rect 150676 3544 150682 3596
rect 156690 3544 156696 3596
rect 156748 3584 156754 3596
rect 164878 3584 164884 3596
rect 156748 3556 164884 3584
rect 156748 3544 156754 3556
rect 164878 3544 164884 3556
rect 164936 3544 164942 3596
rect 173250 3544 173256 3596
rect 173308 3584 173314 3596
rect 475746 3584 475752 3596
rect 173308 3556 475752 3584
rect 173308 3544 173314 3556
rect 475746 3544 475752 3556
rect 475804 3544 475810 3596
rect 508498 3544 508504 3596
rect 508556 3584 508562 3596
rect 524230 3584 524236 3596
rect 508556 3556 524236 3584
rect 508556 3544 508562 3556
rect 524230 3544 524236 3556
rect 524288 3544 524294 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 116670 3516 116676 3528
rect 1728 3488 116676 3516
rect 1728 3476 1734 3488
rect 116670 3476 116676 3488
rect 116728 3476 116734 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 128998 3516 129004 3528
rect 125928 3488 129004 3516
rect 125928 3476 125934 3488
rect 128998 3476 129004 3488
rect 129056 3476 129062 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130654 3516 130660 3528
rect 129424 3488 130660 3516
rect 129424 3476 129430 3488
rect 130654 3476 130660 3488
rect 130712 3476 130718 3528
rect 134702 3476 134708 3528
rect 134760 3516 134766 3528
rect 135254 3516 135260 3528
rect 134760 3488 135260 3516
rect 134760 3476 134766 3488
rect 135254 3476 135260 3488
rect 135312 3476 135318 3528
rect 136266 3476 136272 3528
rect 136324 3516 136330 3528
rect 154206 3516 154212 3528
rect 136324 3488 154212 3516
rect 136324 3476 136330 3488
rect 154206 3476 154212 3488
rect 154264 3476 154270 3528
rect 155218 3476 155224 3528
rect 155276 3516 155282 3528
rect 157794 3516 157800 3528
rect 155276 3488 157800 3516
rect 155276 3476 155282 3488
rect 157794 3476 157800 3488
rect 157852 3476 157858 3528
rect 162118 3476 162124 3528
rect 162176 3516 162182 3528
rect 163682 3516 163688 3528
rect 162176 3488 163688 3516
rect 162176 3476 162182 3488
rect 163682 3476 163688 3488
rect 163740 3476 163746 3528
rect 170582 3476 170588 3528
rect 170640 3516 170646 3528
rect 508866 3516 508872 3528
rect 170640 3488 508872 3516
rect 170640 3476 170646 3488
rect 508866 3476 508872 3488
rect 508924 3476 508930 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 117958 3448 117964 3460
rect 624 3420 117964 3448
rect 624 3408 630 3420
rect 117958 3408 117964 3420
rect 118016 3408 118022 3460
rect 119890 3408 119896 3460
rect 119948 3448 119954 3460
rect 126238 3448 126244 3460
rect 119948 3420 126244 3448
rect 119948 3408 119954 3420
rect 126238 3408 126244 3420
rect 126296 3408 126302 3460
rect 126974 3408 126980 3460
rect 127032 3448 127038 3460
rect 130470 3448 130476 3460
rect 127032 3420 130476 3448
rect 127032 3408 127038 3420
rect 130470 3408 130476 3420
rect 130528 3408 130534 3460
rect 130562 3408 130568 3460
rect 130620 3448 130626 3460
rect 131942 3448 131948 3460
rect 130620 3420 131948 3448
rect 130620 3408 130626 3420
rect 131942 3408 131948 3420
rect 132000 3408 132006 3460
rect 133138 3408 133144 3460
rect 133196 3448 133202 3460
rect 136450 3448 136456 3460
rect 133196 3420 136456 3448
rect 133196 3408 133202 3420
rect 136450 3408 136456 3420
rect 136508 3408 136514 3460
rect 166074 3448 166080 3460
rect 142126 3420 166080 3448
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 18598 3380 18604 3392
rect 17092 3352 18604 3380
rect 17092 3340 17098 3352
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 37182 3340 37188 3392
rect 37240 3380 37246 3392
rect 37918 3380 37924 3392
rect 37240 3352 37924 3380
rect 37240 3340 37246 3352
rect 37918 3340 37924 3352
rect 37976 3340 37982 3392
rect 69106 3340 69112 3392
rect 69164 3380 69170 3392
rect 71038 3380 71044 3392
rect 69164 3352 71044 3380
rect 69164 3340 69170 3352
rect 71038 3340 71044 3352
rect 71096 3340 71102 3392
rect 110506 3340 110512 3392
rect 110564 3380 110570 3392
rect 112438 3380 112444 3392
rect 110564 3352 112444 3380
rect 110564 3340 110570 3352
rect 112438 3340 112444 3352
rect 112496 3340 112502 3392
rect 134058 3340 134064 3392
rect 134116 3380 134122 3392
rect 142126 3380 142154 3420
rect 166074 3408 166080 3420
rect 166132 3408 166138 3460
rect 170490 3408 170496 3460
rect 170548 3448 170554 3460
rect 583386 3448 583392 3460
rect 170548 3420 583392 3448
rect 170548 3408 170554 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 134116 3352 142154 3380
rect 134116 3340 134122 3352
rect 184198 3340 184204 3392
rect 184256 3380 184262 3392
rect 229830 3380 229836 3392
rect 184256 3352 229836 3380
rect 184256 3340 184262 3352
rect 229830 3340 229836 3352
rect 229888 3340 229894 3392
rect 153838 3272 153844 3324
rect 153896 3312 153902 3324
rect 158898 3312 158904 3324
rect 153896 3284 158904 3312
rect 153896 3272 153902 3284
rect 158898 3272 158904 3284
rect 158956 3272 158962 3324
rect 577498 3272 577504 3324
rect 577556 3312 577562 3324
rect 582190 3312 582196 3324
rect 577556 3284 582196 3312
rect 577556 3272 577562 3284
rect 582190 3272 582196 3284
rect 582248 3272 582254 3324
rect 104526 3204 104532 3256
rect 104584 3244 104590 3256
rect 105538 3244 105544 3256
rect 104584 3216 105544 3244
rect 104584 3204 104590 3216
rect 105538 3204 105544 3216
rect 105596 3204 105602 3256
rect 111610 3204 111616 3256
rect 111668 3244 111674 3256
rect 113818 3244 113824 3256
rect 111668 3216 113824 3244
rect 111668 3204 111674 3216
rect 113818 3204 113824 3216
rect 113876 3204 113882 3256
rect 39574 3068 39580 3120
rect 39632 3108 39638 3120
rect 40770 3108 40776 3120
rect 39632 3080 40776 3108
rect 39632 3068 39638 3080
rect 40770 3068 40776 3080
rect 40828 3068 40834 3120
rect 178678 3068 178684 3120
rect 178736 3108 178742 3120
rect 182542 3108 182548 3120
rect 178736 3080 182548 3108
rect 178736 3068 178742 3080
rect 182542 3068 182548 3080
rect 182600 3068 182606 3120
rect 27706 2932 27712 2984
rect 27764 2972 27770 2984
rect 29638 2972 29644 2984
rect 27764 2944 29644 2972
rect 27764 2932 27770 2944
rect 29638 2932 29644 2944
rect 29696 2932 29702 2984
rect 124674 2932 124680 2984
rect 124732 2972 124738 2984
rect 130378 2972 130384 2984
rect 124732 2944 130384 2972
rect 124732 2932 124738 2944
rect 130378 2932 130384 2944
rect 130436 2932 130442 2984
rect 136358 2932 136364 2984
rect 136416 2972 136422 2984
rect 141234 2972 141240 2984
rect 136416 2944 141240 2972
rect 136416 2932 136422 2944
rect 141234 2932 141240 2944
rect 141292 2932 141298 2984
rect 158070 2932 158076 2984
rect 158128 2972 158134 2984
rect 160094 2972 160100 2984
rect 158128 2944 160100 2972
rect 158128 2932 158134 2944
rect 160094 2932 160100 2944
rect 160152 2932 160158 2984
<< via1 >>
rect 332508 700272 332560 700324
rect 397552 700272 397604 700324
rect 194692 700000 194744 700052
rect 202788 700000 202840 700052
rect 260104 699660 260156 699712
rect 267648 699660 267700 699712
rect 193128 696940 193180 696992
rect 194692 696940 194744 696992
rect 188344 694152 188396 694204
rect 193128 694152 193180 694204
rect 253940 690276 253992 690328
rect 260104 690276 260156 690328
rect 238760 683748 238812 683800
rect 253940 683748 253992 683800
rect 233884 679872 233936 679924
rect 238760 679872 238812 679924
rect 183192 679056 183244 679108
rect 188344 679056 188396 679108
rect 180064 677152 180116 677204
rect 183192 677152 183244 677204
rect 175924 657160 175976 657212
rect 180064 657160 180116 657212
rect 156604 643696 156656 643748
rect 175924 643696 175976 643748
rect 150440 635468 150492 635520
rect 156604 635468 156656 635520
rect 141424 631320 141476 631372
rect 150440 631320 150492 631372
rect 3240 605820 3292 605872
rect 43444 605820 43496 605872
rect 211804 591268 211856 591320
rect 233884 591268 233936 591320
rect 422944 590656 422996 590708
rect 579712 590656 579764 590708
rect 209044 580932 209096 580984
rect 211804 580932 211856 580984
rect 134800 574064 134852 574116
rect 141424 574064 141476 574116
rect 127624 570936 127676 570988
rect 134800 570936 134852 570988
rect 195244 570596 195296 570648
rect 209044 570596 209096 570648
rect 189724 567808 189776 567860
rect 195244 567808 195296 567860
rect 3332 553392 3384 553444
rect 43536 553392 43588 553444
rect 124864 552644 124916 552696
rect 127624 552644 127676 552696
rect 396724 536800 396776 536852
rect 580172 536800 580224 536852
rect 119344 532040 119396 532092
rect 124864 532040 124916 532092
rect 184388 511912 184440 511964
rect 189724 511912 189776 511964
rect 114560 511164 114612 511216
rect 119344 511164 119396 511216
rect 117964 508512 118016 508564
rect 137836 508512 137888 508564
rect 178684 507084 178736 507136
rect 184388 507084 184440 507136
rect 112444 504160 112496 504212
rect 114560 504160 114612 504212
rect 116584 487160 116636 487212
rect 117964 487160 118016 487212
rect 418804 484372 418856 484424
rect 580172 484372 580224 484424
rect 174544 482944 174596 482996
rect 178684 482944 178736 482996
rect 115204 472948 115256 473000
rect 116584 472948 116636 473000
rect 166264 467100 166316 467152
rect 174544 467100 174596 467152
rect 93124 461592 93176 461644
rect 112444 461592 112496 461644
rect 162860 452820 162912 452872
rect 166264 452820 166316 452872
rect 2780 449488 2832 449540
rect 4896 449488 4948 449540
rect 155224 447040 155276 447092
rect 162860 447040 162912 447092
rect 442264 444388 442316 444440
rect 580172 444388 580224 444440
rect 79324 436704 79376 436756
rect 93124 436704 93176 436756
rect 413284 430584 413336 430636
rect 580172 430584 580224 430636
rect 76932 419500 76984 419552
rect 79324 419500 79376 419552
rect 73160 417800 73212 417852
rect 76932 417800 76984 417852
rect 64144 413244 64196 413296
rect 73160 413244 73212 413296
rect 152464 411272 152516 411324
rect 155224 411272 155276 411324
rect 50988 404948 51040 405000
rect 64144 404948 64196 405000
rect 47584 401616 47636 401668
rect 50988 401616 51040 401668
rect 3332 397468 3384 397520
rect 13084 397468 13136 397520
rect 46204 382236 46256 382288
rect 47584 382236 47636 382288
rect 421564 378156 421616 378208
rect 580172 378156 580224 378208
rect 115296 363604 115348 363656
rect 152464 363604 152516 363656
rect 58624 356668 58676 356720
rect 115204 356668 115256 356720
rect 45192 350072 45244 350124
rect 46204 350072 46256 350124
rect 2780 345176 2832 345228
rect 5080 345176 5132 345228
rect 57244 339668 57296 339720
rect 58624 339668 58676 339720
rect 95240 337356 95292 337408
rect 115296 337356 115348 337408
rect 93124 328856 93176 328908
rect 95240 328856 95292 328908
rect 55956 327020 56008 327072
rect 57244 327020 57296 327072
rect 417424 324300 417476 324352
rect 579620 324300 579672 324352
rect 54484 321104 54536 321156
rect 55956 321104 56008 321156
rect 53104 309068 53156 309120
rect 54484 309068 54536 309120
rect 87604 304988 87656 305040
rect 93124 304988 93176 305040
rect 3332 292544 3384 292596
rect 43628 292544 43680 292596
rect 73160 287648 73212 287700
rect 87604 287648 87656 287700
rect 57888 280780 57940 280832
rect 73160 280780 73212 280832
rect 51080 279420 51132 279472
rect 53104 279420 53156 279472
rect 47584 277992 47636 278044
rect 57888 277992 57940 278044
rect 48964 273232 49016 273284
rect 50988 273232 51040 273284
rect 410524 271872 410576 271924
rect 579620 271872 579672 271924
rect 46204 270172 46256 270224
rect 47584 270172 47636 270224
rect 47676 262216 47728 262268
rect 48964 262216 49016 262268
rect 46296 259224 46348 259276
rect 47676 259224 47728 259276
rect 45284 249772 45336 249824
rect 46296 249772 46348 249824
rect 3332 240116 3384 240168
rect 21364 240116 21416 240168
rect 44824 225972 44876 226024
rect 72976 225972 73028 226024
rect 45008 224952 45060 225004
rect 68928 224952 68980 225004
rect 45468 224000 45520 224052
rect 46204 224000 46256 224052
rect 45284 215908 45336 215960
rect 56692 215908 56744 215960
rect 57336 215908 57388 215960
rect 68284 215908 68336 215960
rect 45192 214548 45244 214600
rect 57796 214276 57848 214328
rect 174544 211080 174596 211132
rect 176660 211080 176712 211132
rect 177304 210400 177356 210452
rect 580356 210400 580408 210452
rect 45468 209924 45520 209976
rect 47584 209924 47636 209976
rect 57796 209040 57848 209092
rect 69664 209040 69716 209092
rect 68284 208904 68336 208956
rect 75552 208904 75604 208956
rect 69664 204892 69716 204944
rect 85120 204892 85172 204944
rect 47584 202784 47636 202836
rect 51724 202784 51776 202836
rect 75552 201492 75604 201544
rect 78036 201424 78088 201476
rect 85120 201424 85172 201476
rect 87604 201424 87656 201476
rect 78036 198704 78088 198756
rect 81440 198636 81492 198688
rect 81440 194556 81492 194608
rect 84844 194488 84896 194540
rect 87604 194488 87656 194540
rect 89720 194488 89772 194540
rect 89720 191088 89772 191140
rect 111064 191088 111116 191140
rect 149520 191088 149572 191140
rect 266360 191088 266412 191140
rect 147588 189728 147640 189780
rect 236000 189728 236052 189780
rect 146208 188300 146260 188352
rect 207020 188300 207072 188352
rect 3148 187688 3200 187740
rect 112444 187688 112496 187740
rect 144736 185580 144788 185632
rect 174544 185580 174596 185632
rect 84844 184832 84896 184884
rect 86224 184832 86276 184884
rect 134524 183948 134576 184000
rect 137284 183948 137336 184000
rect 111064 182724 111116 182776
rect 113548 182724 113600 182776
rect 151544 182452 151596 182504
rect 154488 182452 154540 182504
rect 138572 182384 138624 182436
rect 154672 182384 154724 182436
rect 133236 181976 133288 182028
rect 136640 181976 136692 182028
rect 146024 181568 146076 181620
rect 136548 181500 136600 181552
rect 118608 181160 118660 181212
rect 138020 181160 138072 181212
rect 113824 181092 113876 181144
rect 137836 181092 137888 181144
rect 137928 181092 137980 181144
rect 138020 181024 138072 181076
rect 128268 180956 128320 181008
rect 146024 180820 146076 180872
rect 113548 180684 113600 180736
rect 116584 180684 116636 180736
rect 146024 180548 146076 180600
rect 155500 180480 155552 180532
rect 161480 180480 161532 180532
rect 155776 180412 155828 180464
rect 163504 180412 163556 180464
rect 155408 180344 155460 180396
rect 163596 180344 163648 180396
rect 129648 179460 129700 179512
rect 136364 179460 136416 179512
rect 86224 179392 86276 179444
rect 133236 179392 133288 179444
rect 140964 179392 141016 179444
rect 89444 179324 89496 179376
rect 120724 178644 120776 178696
rect 136548 178644 136600 178696
rect 162768 177828 162820 177880
rect 164884 177828 164936 177880
rect 154672 177760 154724 177812
rect 121368 177284 121420 177336
rect 137928 177284 137980 177336
rect 141516 177012 141568 177064
rect 146300 177012 146352 177064
rect 161480 176468 161532 176520
rect 124864 175856 124916 175908
rect 138572 175856 138624 175908
rect 161480 175856 161532 175908
rect 161388 174972 161440 175024
rect 161388 174700 161440 174752
rect 89444 173816 89496 173868
rect 92480 173816 92532 173868
rect 161480 167560 161532 167612
rect 161480 167288 161532 167340
rect 92480 167016 92532 167068
rect 95884 166948 95936 167000
rect 51724 164840 51776 164892
rect 66904 164840 66956 164892
rect 147496 162596 147548 162648
rect 136456 161440 136508 161492
rect 137836 161440 137888 161492
rect 161480 161712 161532 161764
rect 163228 161576 163280 161628
rect 164240 161576 164292 161628
rect 160468 161440 160520 161492
rect 161480 161440 161532 161492
rect 135444 161168 135496 161220
rect 136456 161168 136508 161220
rect 163320 159332 163372 159384
rect 173900 159332 173952 159384
rect 133788 158720 133840 158772
rect 136640 158720 136692 158772
rect 132408 158040 132460 158092
rect 135628 158040 135680 158092
rect 131028 157360 131080 157412
rect 134524 157360 134576 157412
rect 136548 157360 136600 157412
rect 138664 157360 138716 157412
rect 151360 157360 151412 157412
rect 152464 157360 152516 157412
rect 66904 155864 66956 155916
rect 69296 155864 69348 155916
rect 95884 155864 95936 155916
rect 97264 155864 97316 155916
rect 148508 155728 148560 155780
rect 148968 155728 149020 155780
rect 69296 152464 69348 152516
rect 84200 152464 84252 152516
rect 84200 149064 84252 149116
rect 87604 149064 87656 149116
rect 164884 146208 164936 146260
rect 165896 146208 165948 146260
rect 124036 137912 124088 137964
rect 124864 137912 124916 137964
rect 146208 137912 146260 137964
rect 147496 137912 147548 137964
rect 152464 137912 152516 137964
rect 155316 137912 155368 137964
rect 134984 137844 135036 137896
rect 136456 137844 136508 137896
rect 150348 137844 150400 137896
rect 153752 137844 153804 137896
rect 148876 137776 148928 137828
rect 152188 137776 152240 137828
rect 156880 137640 156932 137692
rect 163596 137640 163648 137692
rect 161388 137300 161440 137352
rect 170956 137300 171008 137352
rect 162768 137232 162820 137284
rect 172520 137232 172572 137284
rect 158444 137096 158496 137148
rect 163504 137096 163556 137148
rect 119344 136960 119396 137012
rect 120724 136960 120776 137012
rect 148968 136960 149020 137012
rect 150624 136960 150676 137012
rect 147588 136756 147640 136808
rect 149060 136756 149112 136808
rect 160008 136688 160060 136740
rect 161480 136688 161532 136740
rect 3332 136620 3384 136672
rect 112536 136620 112588 136672
rect 45008 135872 45060 135924
rect 178132 135872 178184 135924
rect 116492 129820 116544 129872
rect 116676 129820 116728 129872
rect 97264 129072 97316 129124
rect 102784 129072 102836 129124
rect 102784 117308 102836 117360
rect 105544 117240 105596 117292
rect 87604 104796 87656 104848
rect 90364 104796 90416 104848
rect 116492 100308 116544 100360
rect 116768 100308 116820 100360
rect 90364 99968 90416 100020
rect 101404 99968 101456 100020
rect 177396 99356 177448 99408
rect 580172 99356 580224 99408
rect 105544 92488 105596 92540
rect 109408 92488 109460 92540
rect 109408 89700 109460 89752
rect 101404 89632 101456 89684
rect 104164 89632 104216 89684
rect 114376 89632 114428 89684
rect 3332 84192 3384 84244
rect 116676 84192 116728 84244
rect 175280 76508 175332 76560
rect 527180 76508 527232 76560
rect 43628 75692 43680 75744
rect 114560 75624 114612 75676
rect 119988 75624 120040 75676
rect 13084 75556 13136 75608
rect 4896 75488 4948 75540
rect 135444 74740 135496 74792
rect 421564 75828 421616 75880
rect 170496 75624 170548 75676
rect 170588 75624 170640 75676
rect 170680 75624 170732 75676
rect 177396 75624 177448 75676
rect 170404 75488 170456 75540
rect 170680 75284 170732 75336
rect 417424 75760 417476 75812
rect 135444 74536 135496 74588
rect 143724 74876 143776 74928
rect 146484 74876 146536 74928
rect 143724 74740 143776 74792
rect 172428 75216 172480 75268
rect 462320 75216 462372 75268
rect 170680 74944 170732 74996
rect 170956 74944 171008 74996
rect 580264 75148 580316 75200
rect 168380 74876 168432 74928
rect 172428 74876 172480 74928
rect 157708 74740 157760 74792
rect 169576 74808 169628 74860
rect 169760 74808 169812 74860
rect 170496 74808 170548 74860
rect 170680 74808 170732 74860
rect 235816 74808 235868 74860
rect 249984 74740 250036 74792
rect 285404 74672 285456 74724
rect 112536 74332 112588 74384
rect 148232 74400 148284 74452
rect 116676 74264 116728 74316
rect 148232 74264 148284 74316
rect 112444 74196 112496 74248
rect 152280 74128 152332 74180
rect 152740 74128 152792 74180
rect 148232 74060 148284 74112
rect 139584 73924 139636 73976
rect 141424 73924 141476 73976
rect 140780 73788 140832 73840
rect 141424 73788 141476 73840
rect 152740 73924 152792 73976
rect 153108 73924 153160 73976
rect 320916 74604 320968 74656
rect 343364 74536 343416 74588
rect 167736 74468 167788 74520
rect 413284 74468 413336 74520
rect 167460 74400 167512 74452
rect 410524 74400 410576 74452
rect 170036 74332 170088 74384
rect 169944 74264 169996 74316
rect 168472 74196 168524 74248
rect 397460 74196 397512 74248
rect 159180 74128 159232 74180
rect 484032 74128 484084 74180
rect 170128 74060 170180 74112
rect 171784 74060 171836 74112
rect 515956 74060 516008 74112
rect 163044 73992 163096 74044
rect 533712 73992 533764 74044
rect 164424 73924 164476 73976
rect 551468 73924 551520 73976
rect 163320 73856 163372 73908
rect 537208 73856 537260 73908
rect 164700 73788 164752 73840
rect 554964 73788 555016 73840
rect 5080 73720 5132 73772
rect 140964 73652 141016 73704
rect 161664 73720 161716 73772
rect 171784 73720 171836 73772
rect 140780 73584 140832 73636
rect 141056 73584 141108 73636
rect 141700 73584 141752 73636
rect 140964 73448 141016 73500
rect 141240 73448 141292 73500
rect 141148 73380 141200 73432
rect 141516 73380 141568 73432
rect 122932 73312 122984 73364
rect 123668 73312 123720 73364
rect 141240 73312 141292 73364
rect 169668 73652 169720 73704
rect 167920 73584 167972 73636
rect 172704 73584 172756 73636
rect 167644 73516 167696 73568
rect 170588 73516 170640 73568
rect 168104 73448 168156 73500
rect 170956 73448 171008 73500
rect 142068 73380 142120 73432
rect 158904 73312 158956 73364
rect 163044 73312 163096 73364
rect 124312 73176 124364 73228
rect 113916 72768 113968 72820
rect 141424 73108 141476 73160
rect 142344 73108 142396 73160
rect 143080 73108 143132 73160
rect 150440 73176 150492 73228
rect 119620 73040 119672 73092
rect 130384 73040 130436 73092
rect 147772 73040 147824 73092
rect 148232 73040 148284 73092
rect 121184 72972 121236 73024
rect 129280 72972 129332 73024
rect 136640 72972 136692 73024
rect 139860 72972 139912 73024
rect 123116 72904 123168 72956
rect 123576 72904 123628 72956
rect 121276 72768 121328 72820
rect 125232 72836 125284 72888
rect 129740 72904 129792 72956
rect 129924 72904 129976 72956
rect 130384 72904 130436 72956
rect 130568 72904 130620 72956
rect 129832 72836 129884 72888
rect 145104 72836 145156 72888
rect 130292 72768 130344 72820
rect 130568 72768 130620 72820
rect 118148 72700 118200 72752
rect 123760 72700 123812 72752
rect 124588 72700 124640 72752
rect 125232 72700 125284 72752
rect 125508 72700 125560 72752
rect 126428 72700 126480 72752
rect 126796 72700 126848 72752
rect 129924 72700 129976 72752
rect 130108 72700 130160 72752
rect 134616 72700 134668 72752
rect 135076 72700 135128 72752
rect 145104 72700 145156 72752
rect 145840 72700 145892 72752
rect 109684 72632 109736 72684
rect 107016 72496 107068 72548
rect 123024 72496 123076 72548
rect 123392 72632 123444 72684
rect 123208 72564 123260 72616
rect 124864 72632 124916 72684
rect 141608 72632 141660 72684
rect 141792 72632 141844 72684
rect 152280 73244 152332 73296
rect 151360 73176 151412 73228
rect 152280 73108 152332 73160
rect 153292 73108 153344 73160
rect 152372 72972 152424 73024
rect 153108 72836 153160 72888
rect 152372 72768 152424 72820
rect 152648 72768 152700 72820
rect 151084 72700 151136 72752
rect 151360 72700 151412 72752
rect 151636 72700 151688 72752
rect 158812 73244 158864 73296
rect 157984 73176 158036 73228
rect 154948 73108 155000 73160
rect 157708 73108 157760 73160
rect 158812 73108 158864 73160
rect 168380 73244 168432 73296
rect 168840 73244 168892 73296
rect 160836 73176 160888 73228
rect 505376 73176 505428 73228
rect 164424 73108 164476 73160
rect 168288 73108 168340 73160
rect 175280 73108 175332 73160
rect 155500 73040 155552 73092
rect 156052 73040 156104 73092
rect 158904 73040 158956 73092
rect 159180 73040 159232 73092
rect 160008 73040 160060 73092
rect 165712 73040 165764 73092
rect 166908 73040 166960 73092
rect 167828 73040 167880 73092
rect 178684 73040 178736 73092
rect 153844 72768 153896 72820
rect 155500 72768 155552 72820
rect 167552 72972 167604 73024
rect 168012 72972 168064 73024
rect 172152 72972 172204 73024
rect 172336 72972 172388 73024
rect 157156 72904 157208 72956
rect 168932 72904 168984 72956
rect 422944 72972 422996 73024
rect 178684 72904 178736 72956
rect 418804 72904 418856 72956
rect 162584 72836 162636 72888
rect 157524 72768 157576 72820
rect 159456 72768 159508 72820
rect 160008 72768 160060 72820
rect 160284 72768 160336 72820
rect 160744 72768 160796 72820
rect 172704 72836 172756 72888
rect 396724 72836 396776 72888
rect 167736 72768 167788 72820
rect 168472 72768 168524 72820
rect 168748 72768 168800 72820
rect 162584 72700 162636 72752
rect 168104 72700 168156 72752
rect 168564 72700 168616 72752
rect 397552 72768 397604 72820
rect 167644 72632 167696 72684
rect 168196 72632 168248 72684
rect 177304 72632 177356 72684
rect 123576 72564 123628 72616
rect 150440 72564 150492 72616
rect 152648 72564 152700 72616
rect 152924 72564 152976 72616
rect 153108 72564 153160 72616
rect 124312 72496 124364 72548
rect 153844 72496 153896 72548
rect 154672 72564 154724 72616
rect 154856 72564 154908 72616
rect 156144 72564 156196 72616
rect 445024 72564 445076 72616
rect 161848 72496 161900 72548
rect 162584 72496 162636 72548
rect 163412 72496 163464 72548
rect 163596 72496 163648 72548
rect 164424 72496 164476 72548
rect 471244 72496 471296 72548
rect 23020 72428 23072 72480
rect 123300 72428 123352 72480
rect 123392 72428 123444 72480
rect 153292 72428 153344 72480
rect 157248 72428 157300 72480
rect 160836 72428 160888 72480
rect 161388 72428 161440 72480
rect 161940 72428 161992 72480
rect 162676 72428 162728 72480
rect 163136 72428 163188 72480
rect 163964 72428 164016 72480
rect 166816 72428 166868 72480
rect 580264 72428 580316 72480
rect 121000 72292 121052 72344
rect 127900 72360 127952 72412
rect 130108 72360 130160 72412
rect 130660 72360 130712 72412
rect 133052 72360 133104 72412
rect 133604 72360 133656 72412
rect 148232 72360 148284 72412
rect 148600 72360 148652 72412
rect 152188 72360 152240 72412
rect 123392 72292 123444 72344
rect 124128 72292 124180 72344
rect 120908 72224 120960 72276
rect 128176 72292 128228 72344
rect 132592 72292 132644 72344
rect 133512 72292 133564 72344
rect 135904 72292 135956 72344
rect 136272 72292 136324 72344
rect 149704 72292 149756 72344
rect 153292 72292 153344 72344
rect 124404 72224 124456 72276
rect 126244 72224 126296 72276
rect 150256 72224 150308 72276
rect 152188 72224 152240 72276
rect 124128 72156 124180 72208
rect 126704 72156 126756 72208
rect 127440 72156 127492 72208
rect 127808 72156 127860 72208
rect 149152 72156 149204 72208
rect 154488 72156 154540 72208
rect 123576 72088 123628 72140
rect 125968 72088 126020 72140
rect 135444 72088 135496 72140
rect 135628 72088 135680 72140
rect 138112 72088 138164 72140
rect 139308 72088 139360 72140
rect 157708 72360 157760 72412
rect 168196 72360 168248 72412
rect 156604 72292 156656 72344
rect 169116 72292 169168 72344
rect 156144 72224 156196 72276
rect 158628 72224 158680 72276
rect 160928 72224 160980 72276
rect 161204 72224 161256 72276
rect 155500 72156 155552 72208
rect 161940 72156 161992 72208
rect 163044 72156 163096 72208
rect 169208 72156 169260 72208
rect 158260 72088 158312 72140
rect 167368 72088 167420 72140
rect 580816 72088 580868 72140
rect 119344 72020 119396 72072
rect 129740 72020 129792 72072
rect 132684 72020 132736 72072
rect 134524 72020 134576 72072
rect 160376 72020 160428 72072
rect 160928 72020 160980 72072
rect 164608 72020 164660 72072
rect 165160 72020 165212 72072
rect 167000 72020 167052 72072
rect 580172 72020 580224 72072
rect 122840 71952 122892 72004
rect 131120 71952 131172 72004
rect 154396 71952 154448 72004
rect 167920 71952 167972 72004
rect 120724 71884 120776 71936
rect 126980 71884 127032 71936
rect 151912 71884 151964 71936
rect 116768 71816 116820 71868
rect 123208 71816 123260 71868
rect 127716 71816 127768 71868
rect 131028 71816 131080 71868
rect 149060 71816 149112 71868
rect 118056 71748 118108 71800
rect 122932 71748 122984 71800
rect 128176 71748 128228 71800
rect 131488 71748 131540 71800
rect 146024 71748 146076 71800
rect 149704 71748 149756 71800
rect 156328 71748 156380 71800
rect 156880 71748 156932 71800
rect 158904 71884 158956 71936
rect 168012 71884 168064 71936
rect 157524 71816 157576 71868
rect 161940 71816 161992 71868
rect 167828 71816 167880 71868
rect 157708 71748 157760 71800
rect 158904 71748 158956 71800
rect 160744 71748 160796 71800
rect 165620 71748 165672 71800
rect 119436 71680 119488 71732
rect 122748 71680 122800 71732
rect 155500 71680 155552 71732
rect 165712 71680 165764 71732
rect 171784 71680 171836 71732
rect 171876 71680 171928 71732
rect 580448 71680 580500 71732
rect 120816 71612 120868 71664
rect 126428 71612 126480 71664
rect 140780 71612 140832 71664
rect 251180 71612 251232 71664
rect 117964 71544 118016 71596
rect 124772 71544 124824 71596
rect 140964 71544 141016 71596
rect 253480 71544 253532 71596
rect 143540 71476 143592 71528
rect 283104 71476 283156 71528
rect 144000 71408 144052 71460
rect 288992 71408 289044 71460
rect 145472 71340 145524 71392
rect 307944 71340 307996 71392
rect 121092 71272 121144 71324
rect 130936 71272 130988 71324
rect 152004 71272 152056 71324
rect 391848 71272 391900 71324
rect 111064 71204 111116 71256
rect 129188 71204 129240 71256
rect 84476 71136 84528 71188
rect 128084 71136 128136 71188
rect 156420 71136 156472 71188
rect 448612 71204 448664 71256
rect 161388 71136 161440 71188
rect 504180 71136 504232 71188
rect 41880 71068 41932 71120
rect 117964 71068 118016 71120
rect 167736 71068 167788 71120
rect 168196 71068 168248 71120
rect 171784 71068 171836 71120
rect 538404 71068 538456 71120
rect 29644 71000 29696 71052
rect 142344 71000 142396 71052
rect 139860 70932 139912 70984
rect 164148 71000 164200 71052
rect 545488 71000 545540 71052
rect 123760 70864 123812 70916
rect 145564 70864 145616 70916
rect 145840 70864 145892 70916
rect 247592 70932 247644 70984
rect 194416 70864 194468 70916
rect 136088 70796 136140 70848
rect 170404 70796 170456 70848
rect 116400 70728 116452 70780
rect 130384 70728 130436 70780
rect 167092 70728 167144 70780
rect 171876 70728 171928 70780
rect 157984 70660 158036 70712
rect 167736 70660 167788 70712
rect 130384 70456 130436 70508
rect 131212 70456 131264 70508
rect 121736 70388 121788 70440
rect 122104 70388 122156 70440
rect 3516 70320 3568 70372
rect 169392 70320 169444 70372
rect 43536 70252 43588 70304
rect 162216 70252 162268 70304
rect 145748 70184 145800 70236
rect 311440 70184 311492 70236
rect 134708 70116 134760 70168
rect 118792 69980 118844 70032
rect 130752 69980 130804 70032
rect 80888 69844 80940 69896
rect 127440 69844 127492 69896
rect 71044 69776 71096 69828
rect 126888 69776 126940 69828
rect 54944 69708 54996 69760
rect 125784 69708 125836 69760
rect 47860 69640 47912 69692
rect 124220 69640 124272 69692
rect 155500 70116 155552 70168
rect 354036 70116 354088 70168
rect 151268 70048 151320 70100
rect 382372 70048 382424 70100
rect 157248 69980 157300 70032
rect 396540 69980 396592 70032
rect 153200 69912 153252 69964
rect 161940 69912 161992 69964
rect 403624 69912 403676 69964
rect 407212 69844 407264 69896
rect 157800 69776 157852 69828
rect 466276 69776 466328 69828
rect 158076 69708 158128 69760
rect 469864 69708 469916 69760
rect 160192 69640 160244 69692
rect 497096 69640 497148 69692
rect 148508 69572 148560 69624
rect 189816 69572 189868 69624
rect 116584 69436 116636 69488
rect 152648 69164 152700 69216
rect 161940 69164 161992 69216
rect 169576 69300 169628 69352
rect 162216 69232 162268 69284
rect 169300 69232 169352 69284
rect 168472 69164 168524 69216
rect 119528 69028 119580 69080
rect 125232 69028 125284 69080
rect 134616 68824 134668 68876
rect 167184 68824 167236 68876
rect 135444 68756 135496 68808
rect 181444 68756 181496 68808
rect 117596 68688 117648 68740
rect 130108 68688 130160 68740
rect 139308 68688 139360 68740
rect 213368 68688 213420 68740
rect 113824 68620 113876 68672
rect 130200 68620 130252 68672
rect 140320 68620 140372 68672
rect 241704 68620 241756 68672
rect 105544 68552 105596 68604
rect 129648 68552 129700 68604
rect 157432 68552 157484 68604
rect 461584 68552 461636 68604
rect 93952 68484 94004 68536
rect 128820 68484 128872 68536
rect 164700 68484 164752 68536
rect 553768 68484 553820 68536
rect 58440 68416 58492 68468
rect 126060 68416 126112 68468
rect 133144 68416 133196 68468
rect 135904 68416 135956 68468
rect 164608 68416 164660 68468
rect 560852 68416 560904 68468
rect 30104 68348 30156 68400
rect 123852 68348 123904 68400
rect 166908 68348 166960 68400
rect 568028 68348 568080 68400
rect 7656 68280 7708 68332
rect 121736 68280 121788 68332
rect 166264 68280 166316 68332
rect 575112 68280 575164 68332
rect 141056 68076 141108 68128
rect 141516 68076 141568 68128
rect 130476 67600 130528 67652
rect 131396 67600 131448 67652
rect 150808 67532 150860 67584
rect 151544 67532 151596 67584
rect 142804 67464 142856 67516
rect 143080 67464 143132 67516
rect 155960 67464 156012 67516
rect 156788 67464 156840 67516
rect 115204 67124 115256 67176
rect 130292 67124 130344 67176
rect 161296 67124 161348 67176
rect 170588 67124 170640 67176
rect 103336 67056 103388 67108
rect 129556 67056 129608 67108
rect 146944 67056 146996 67108
rect 326804 67056 326856 67108
rect 332600 67056 332652 67108
rect 472256 67056 472308 67108
rect 97448 66988 97500 67040
rect 129096 66988 129148 67040
rect 141240 66988 141292 67040
rect 141700 66988 141752 67040
rect 148876 66988 148928 67040
rect 348056 66988 348108 67040
rect 76196 66920 76248 66972
rect 127072 66920 127124 66972
rect 154488 66920 154540 66972
rect 355232 66920 355284 66972
rect 60832 66852 60884 66904
rect 124404 66852 124456 66904
rect 141700 66852 141752 66904
rect 141884 66852 141936 66904
rect 145564 66852 145616 66904
rect 145932 66852 145984 66904
rect 152188 66852 152240 66904
rect 369400 66852 369452 66904
rect 137100 66716 137152 66768
rect 137744 66716 137796 66768
rect 129188 66240 129240 66292
rect 131304 66240 131356 66292
rect 121920 65968 121972 66020
rect 122196 65968 122248 66020
rect 132868 65968 132920 66020
rect 134616 65968 134668 66020
rect 121552 65900 121604 65952
rect 128268 65900 128320 65952
rect 128820 65900 128872 65952
rect 129004 65900 129056 65952
rect 138756 65900 138808 65952
rect 139216 65900 139268 65952
rect 142712 65900 142764 65952
rect 142988 65900 143040 65952
rect 112444 65832 112496 65884
rect 129924 65832 129976 65884
rect 139952 65832 140004 65884
rect 140412 65832 140464 65884
rect 154948 65832 155000 65884
rect 155776 65832 155828 65884
rect 159732 65832 159784 65884
rect 166908 65832 166960 65884
rect 101036 65764 101088 65816
rect 129372 65764 129424 65816
rect 134248 65764 134300 65816
rect 134892 65764 134944 65816
rect 135076 65764 135128 65816
rect 168380 65764 168432 65816
rect 86868 65696 86920 65748
rect 121552 65696 121604 65748
rect 79692 65628 79744 65680
rect 127900 65696 127952 65748
rect 121828 65628 121880 65680
rect 122380 65628 122432 65680
rect 123300 65628 123352 65680
rect 123944 65628 123996 65680
rect 127532 65628 127584 65680
rect 127808 65628 127860 65680
rect 26516 65560 26568 65612
rect 123116 65560 123168 65612
rect 2872 65492 2924 65544
rect 121644 65492 121696 65544
rect 121736 65492 121788 65544
rect 122564 65492 122616 65544
rect 125140 65492 125192 65544
rect 125508 65492 125560 65544
rect 126152 65492 126204 65544
rect 126612 65492 126664 65544
rect 128728 65492 128780 65544
rect 129280 65492 129332 65544
rect 130660 65492 130712 65544
rect 131580 65492 131632 65544
rect 131948 65492 132000 65544
rect 132316 65492 132368 65544
rect 133420 65696 133472 65748
rect 134340 65696 134392 65748
rect 134800 65696 134852 65748
rect 137100 65696 137152 65748
rect 137652 65696 137704 65748
rect 139768 65696 139820 65748
rect 140320 65696 140372 65748
rect 136824 65628 136876 65680
rect 137468 65628 137520 65680
rect 138388 65628 138440 65680
rect 138572 65628 138624 65680
rect 139400 65628 139452 65680
rect 184204 65696 184256 65748
rect 144000 65628 144052 65680
rect 144276 65628 144328 65680
rect 149336 65628 149388 65680
rect 150164 65628 150216 65680
rect 150532 65628 150584 65680
rect 151268 65628 151320 65680
rect 153568 65628 153620 65680
rect 154396 65628 154448 65680
rect 155132 65628 155184 65680
rect 123484 65356 123536 65408
rect 123852 65356 123904 65408
rect 129004 65356 129056 65408
rect 129188 65356 129240 65408
rect 131856 65356 131908 65408
rect 132132 65356 132184 65408
rect 132592 65356 132644 65408
rect 131764 65288 131816 65340
rect 132776 65560 132828 65612
rect 134064 65560 134116 65612
rect 134432 65560 134484 65612
rect 135628 65560 135680 65612
rect 136180 65560 136232 65612
rect 137284 65560 137336 65612
rect 137652 65560 137704 65612
rect 133972 65492 134024 65544
rect 134984 65492 135036 65544
rect 136916 65492 136968 65544
rect 137468 65492 137520 65544
rect 132776 65356 132828 65408
rect 133420 65356 133472 65408
rect 135352 65356 135404 65408
rect 136088 65356 136140 65408
rect 133420 65220 133472 65272
rect 142252 65560 142304 65612
rect 143264 65560 143316 65612
rect 143632 65560 143684 65612
rect 144552 65560 144604 65612
rect 144920 65560 144972 65612
rect 145748 65560 145800 65612
rect 148048 65560 148100 65612
rect 148784 65560 148836 65612
rect 138940 65492 138992 65544
rect 139124 65492 139176 65544
rect 139492 65492 139544 65544
rect 140504 65492 140556 65544
rect 140872 65492 140924 65544
rect 141792 65492 141844 65544
rect 142436 65492 142488 65544
rect 143172 65492 143224 65544
rect 144092 65492 144144 65544
rect 144644 65492 144696 65544
rect 145196 65492 145248 65544
rect 145840 65492 145892 65544
rect 147680 65492 147732 65544
rect 148140 65492 148192 65544
rect 148324 65492 148376 65544
rect 148692 65492 148744 65544
rect 139860 65424 139912 65476
rect 140228 65424 140280 65476
rect 149888 65560 149940 65612
rect 153200 65560 153252 65612
rect 154028 65560 154080 65612
rect 154672 65560 154724 65612
rect 155224 65560 155276 65612
rect 149612 65492 149664 65544
rect 149980 65492 150032 65544
rect 150532 65492 150584 65544
rect 150992 65492 151044 65544
rect 151820 65492 151872 65544
rect 152924 65492 152976 65544
rect 153752 65492 153804 65544
rect 154212 65492 154264 65544
rect 138940 65356 138992 65408
rect 143908 65356 143960 65408
rect 144368 65356 144420 65408
rect 146668 65356 146720 65408
rect 147220 65356 147272 65408
rect 149428 65356 149480 65408
rect 146852 65288 146904 65340
rect 147312 65288 147364 65340
rect 151176 65424 151228 65476
rect 153476 65424 153528 65476
rect 154304 65424 154356 65476
rect 156236 65628 156288 65680
rect 446220 65628 446272 65680
rect 160100 65560 160152 65612
rect 161112 65560 161164 65612
rect 162032 65560 162084 65612
rect 162492 65560 162544 65612
rect 163228 65560 163280 65612
rect 163688 65560 163740 65612
rect 164240 65560 164292 65612
rect 165252 65560 165304 65612
rect 165620 65560 165672 65612
rect 166724 65560 166776 65612
rect 157432 65492 157484 65544
rect 157892 65492 157944 65544
rect 158720 65492 158772 65544
rect 159180 65492 159232 65544
rect 160468 65492 160520 65544
rect 160836 65492 160888 65544
rect 162860 65492 162912 65544
rect 164056 65492 164108 65544
rect 164516 65492 164568 65544
rect 165068 65492 165120 65544
rect 165804 65492 165856 65544
rect 166540 65492 166592 65544
rect 160008 65424 160060 65476
rect 155408 65356 155460 65408
rect 159272 65356 159324 65408
rect 159732 65356 159784 65408
rect 163412 65356 163464 65408
rect 163872 65356 163924 65408
rect 164332 65424 164384 65476
rect 165344 65424 165396 65476
rect 487620 65560 487672 65612
rect 166908 65492 166960 65544
rect 491116 65492 491168 65544
rect 165712 65356 165764 65408
rect 166264 65356 166316 65408
rect 154856 65288 154908 65340
rect 155592 65288 155644 65340
rect 163320 65288 163372 65340
rect 163780 65288 163832 65340
rect 138664 65220 138716 65272
rect 139032 65220 139084 65272
rect 139584 65220 139636 65272
rect 140320 65220 140372 65272
rect 142528 65220 142580 65272
rect 142896 65220 142948 65272
rect 146300 65220 146352 65272
rect 147128 65220 147180 65272
rect 147864 65220 147916 65272
rect 148324 65220 148376 65272
rect 151084 65220 151136 65272
rect 154580 65220 154632 65272
rect 155500 65220 155552 65272
rect 158904 65220 158956 65272
rect 159364 65220 159416 65272
rect 161664 65220 161716 65272
rect 162216 65220 162268 65272
rect 162952 65220 163004 65272
rect 163872 65220 163924 65272
rect 138756 65152 138808 65204
rect 158996 65152 159048 65204
rect 159548 65152 159600 65204
rect 131764 65084 131816 65136
rect 138020 65084 138072 65136
rect 138848 65084 138900 65136
rect 158812 65084 158864 65136
rect 159456 65084 159508 65136
rect 138204 64948 138256 65000
rect 138940 64948 138992 65000
rect 112812 64336 112864 64388
rect 130568 64336 130620 64388
rect 67916 64268 67968 64320
rect 124128 64268 124180 64320
rect 135720 64268 135772 64320
rect 178684 64268 178736 64320
rect 48964 64200 49016 64252
rect 125324 64200 125376 64252
rect 152372 64200 152424 64252
rect 152464 64200 152516 64252
rect 397736 64200 397788 64252
rect 12348 64132 12400 64184
rect 122472 64132 122524 64184
rect 162676 64132 162728 64184
rect 519544 64132 519596 64184
rect 152372 63996 152424 64048
rect 146392 63724 146444 63776
rect 147036 63724 147088 63776
rect 161848 63452 161900 63504
rect 162400 63452 162452 63504
rect 156420 63316 156472 63368
rect 157064 63316 157116 63368
rect 137744 63044 137796 63096
rect 200304 63044 200356 63096
rect 4804 62976 4856 63028
rect 170312 62976 170364 63028
rect 102232 62908 102284 62960
rect 129464 62908 129516 62960
rect 136732 62908 136784 62960
rect 137744 62908 137796 62960
rect 149060 62908 149112 62960
rect 356336 62908 356388 62960
rect 56048 62840 56100 62892
rect 125876 62840 125928 62892
rect 158260 62840 158312 62892
rect 394240 62840 394292 62892
rect 44272 62772 44324 62824
rect 124956 62772 125008 62824
rect 162768 62772 162820 62824
rect 523040 62772 523092 62824
rect 133236 62024 133288 62076
rect 135996 62024 136048 62076
rect 109316 61480 109368 61532
rect 130016 61480 130068 61532
rect 139216 61480 139268 61532
rect 221556 61480 221608 61532
rect 65524 61412 65576 61464
rect 126704 61412 126756 61464
rect 150624 61412 150676 61464
rect 374092 61412 374144 61464
rect 40684 61344 40736 61396
rect 124680 61344 124732 61396
rect 156696 61344 156748 61396
rect 453304 61344 453356 61396
rect 157708 61140 157760 61192
rect 157984 61140 158036 61192
rect 149796 61072 149848 61124
rect 150072 61072 150124 61124
rect 117228 60800 117280 60852
rect 122288 60800 122340 60852
rect 137192 60188 137244 60240
rect 207388 60188 207440 60240
rect 63224 60120 63276 60172
rect 126796 60120 126848 60172
rect 140136 60120 140188 60172
rect 239312 60120 239364 60172
rect 59636 60052 59688 60104
rect 126612 60052 126664 60104
rect 148324 60052 148376 60104
rect 338672 60052 338724 60104
rect 9956 59984 10008 60036
rect 117228 59984 117280 60036
rect 126244 59984 126296 60036
rect 130844 59984 130896 60036
rect 151084 59984 151136 60036
rect 381176 59984 381228 60036
rect 135260 58896 135312 58948
rect 176660 58896 176712 58948
rect 152464 58828 152516 58880
rect 277124 58828 277176 58880
rect 153936 58760 153988 58812
rect 409604 58760 409656 58812
rect 163412 58692 163464 58744
rect 544384 58692 544436 58744
rect 25320 58624 25372 58676
rect 123852 58624 123904 58676
rect 166448 58624 166500 58676
rect 572720 58624 572772 58676
rect 114008 58352 114060 58404
rect 119620 58352 119672 58404
rect 133236 57876 133288 57928
rect 136364 57876 136416 57928
rect 138664 57400 138716 57452
rect 225144 57400 225196 57452
rect 106924 57332 106976 57384
rect 121276 57332 121328 57384
rect 142712 57332 142764 57384
rect 271236 57332 271288 57384
rect 77392 57264 77444 57316
rect 127808 57264 127860 57316
rect 145564 57264 145616 57316
rect 313832 57264 313884 57316
rect 8760 57196 8812 57248
rect 121828 57196 121880 57248
rect 163504 57196 163556 57248
rect 540796 57196 540848 57248
rect 136088 55972 136140 56024
rect 177856 55972 177908 56024
rect 57244 55904 57296 55956
rect 123576 55904 123628 55956
rect 149612 55904 149664 55956
rect 359924 55904 359976 55956
rect 32404 55836 32456 55888
rect 123760 55836 123812 55888
rect 164976 55836 165028 55888
rect 558552 55836 558604 55888
rect 138756 54748 138808 54800
rect 216864 54748 216916 54800
rect 142804 54680 142856 54732
rect 274824 54680 274876 54732
rect 146852 54612 146904 54664
rect 324412 54612 324464 54664
rect 155132 54544 155184 54596
rect 427268 54544 427320 54596
rect 33600 54476 33652 54528
rect 123392 54476 123444 54528
rect 159456 54476 159508 54528
rect 468668 54476 468720 54528
rect 136180 53456 136232 53508
rect 186136 53456 186188 53508
rect 137284 53388 137336 53440
rect 201500 53388 201552 53440
rect 148416 53320 148468 53372
rect 342168 53320 342220 53372
rect 154028 53252 154080 53304
rect 413100 53252 413152 53304
rect 163596 53184 163648 53236
rect 539600 53184 539652 53236
rect 62028 53116 62080 53168
rect 126336 53116 126388 53168
rect 165068 53116 165120 53168
rect 552664 53116 552716 53168
rect 31300 53048 31352 53100
rect 123300 53048 123352 53100
rect 166540 53048 166592 53100
rect 569132 53048 569184 53100
rect 133328 52436 133380 52488
rect 136180 52436 136232 52488
rect 132040 52368 132092 52420
rect 134708 52368 134760 52420
rect 146944 51892 146996 51944
rect 328000 51892 328052 51944
rect 151176 51824 151228 51876
rect 377680 51824 377732 51876
rect 167552 51756 167604 51808
rect 436744 51756 436796 51808
rect 13544 51688 13596 51740
rect 121736 51688 121788 51740
rect 162124 51688 162176 51740
rect 508504 51688 508556 51740
rect 137376 50600 137428 50652
rect 203892 50600 203944 50652
rect 145656 50532 145708 50584
rect 310244 50532 310296 50584
rect 149796 50464 149848 50516
rect 367008 50464 367060 50516
rect 155224 50396 155276 50448
rect 430856 50396 430908 50448
rect 14740 50328 14792 50380
rect 122656 50328 122708 50380
rect 165160 50328 165212 50380
rect 562048 50328 562100 50380
rect 136272 49036 136324 49088
rect 184940 49036 184992 49088
rect 99840 48968 99892 49020
rect 121184 48968 121236 49020
rect 148508 48968 148560 49020
rect 345756 48968 345808 49020
rect 135444 47812 135496 47864
rect 180248 47812 180300 47864
rect 144184 47744 144236 47796
rect 291384 47744 291436 47796
rect 149888 47676 149940 47728
rect 363512 47676 363564 47728
rect 92756 47608 92808 47660
rect 129280 47608 129332 47660
rect 154120 47608 154172 47660
rect 416688 47608 416740 47660
rect 83280 47540 83332 47592
rect 127992 47540 128044 47592
rect 156788 47540 156840 47592
rect 442632 47540 442684 47592
rect 135628 46248 135680 46300
rect 188528 46248 188580 46300
rect 4068 46180 4120 46232
rect 122288 46180 122340 46232
rect 140228 46180 140280 46232
rect 234620 46180 234672 46232
rect 3424 45500 3476 45552
rect 170220 45500 170272 45552
rect 152740 44956 152792 45008
rect 398932 44956 398984 45008
rect 95148 44888 95200 44940
rect 129096 44888 129148 44940
rect 156880 44888 156932 44940
rect 447416 44888 447468 44940
rect 64328 44820 64380 44872
rect 126520 44820 126572 44872
rect 160836 44820 160888 44872
rect 500592 44820 500644 44872
rect 137468 43596 137520 43648
rect 197912 43596 197964 43648
rect 155316 43528 155368 43580
rect 434444 43528 434496 43580
rect 159548 43460 159600 43512
rect 481732 43460 481784 43512
rect 133420 43392 133472 43444
rect 144736 43392 144788 43444
rect 162216 43392 162268 43444
rect 514760 43392 514812 43444
rect 132132 42712 132184 42764
rect 132960 42712 133012 42764
rect 138848 42236 138900 42288
rect 212172 42236 212224 42288
rect 149980 42168 150032 42220
rect 361120 42168 361172 42220
rect 152832 42100 152884 42152
rect 402520 42100 402572 42152
rect 162308 42032 162360 42084
rect 525432 42032 525484 42084
rect 138940 40876 138992 40928
rect 215668 40876 215720 40928
rect 142896 40808 142948 40860
rect 270040 40808 270092 40860
rect 159640 40740 159692 40792
rect 486424 40740 486476 40792
rect 82084 40672 82136 40724
rect 121000 40672 121052 40724
rect 134432 40672 134484 40724
rect 160744 40672 160796 40724
rect 160928 40672 160980 40724
rect 499396 40672 499448 40724
rect 135812 39516 135864 39568
rect 183744 39516 183796 39568
rect 143816 39448 143868 39500
rect 286600 39448 286652 39500
rect 161020 39380 161072 39432
rect 506480 39380 506532 39432
rect 163688 39312 163740 39364
rect 543188 39312 543240 39364
rect 137560 38088 137612 38140
rect 206192 38088 206244 38140
rect 145748 38020 145800 38072
rect 300768 38020 300820 38072
rect 153844 37952 153896 38004
rect 362316 37952 362368 38004
rect 166632 37884 166684 37936
rect 573916 37884 573968 37936
rect 141424 36660 141476 36712
rect 259460 36660 259512 36712
rect 134800 36592 134852 36644
rect 156696 36592 156748 36644
rect 168288 36592 168340 36644
rect 429660 36592 429712 36644
rect 155408 36524 155460 36576
rect 432052 36524 432104 36576
rect 142988 35368 143040 35420
rect 272432 35368 272484 35420
rect 147036 35300 147088 35352
rect 319720 35300 319772 35352
rect 169208 35232 169260 35284
rect 465172 35232 465224 35284
rect 161112 35164 161164 35216
rect 495900 35164 495952 35216
rect 143080 33872 143132 33924
rect 273628 33872 273680 33924
rect 155500 33804 155552 33856
rect 424968 33804 425020 33856
rect 162400 33736 162452 33788
rect 517152 33736 517204 33788
rect 139032 32648 139084 32700
rect 219256 32648 219308 32700
rect 144276 32580 144328 32632
rect 293684 32580 293736 32632
rect 148600 32512 148652 32564
rect 337476 32512 337528 32564
rect 162584 32444 162636 32496
rect 518348 32444 518400 32496
rect 133512 32376 133564 32428
rect 142436 32376 142488 32428
rect 162492 32376 162544 32428
rect 520740 32376 520792 32428
rect 140320 31288 140372 31340
rect 233424 31288 233476 31340
rect 150072 31220 150124 31272
rect 357532 31220 357584 31272
rect 159732 31152 159784 31204
rect 485228 31152 485280 31204
rect 163780 31084 163832 31136
rect 536104 31084 536156 31136
rect 134892 31016 134944 31068
rect 162124 31016 162176 31068
rect 165252 31016 165304 31068
rect 549076 31016 549128 31068
rect 134984 29724 135036 29776
rect 158076 29724 158128 29776
rect 156972 29656 157024 29708
rect 454500 29656 454552 29708
rect 157340 29588 157392 29640
rect 460388 29588 460440 29640
rect 139124 28568 139176 28620
rect 223948 28568 224000 28620
rect 143172 28500 143224 28552
rect 268844 28500 268896 28552
rect 151268 28432 151320 28484
rect 372896 28432 372948 28484
rect 155960 28364 156012 28416
rect 449808 28364 449860 28416
rect 159824 28296 159876 28348
rect 488816 28296 488868 28348
rect 166724 28228 166776 28280
rect 566832 28228 566884 28280
rect 149704 27072 149756 27124
rect 315028 27072 315080 27124
rect 151360 27004 151412 27056
rect 379980 27004 380032 27056
rect 160376 26936 160428 26988
rect 507676 26936 507728 26988
rect 165896 26868 165948 26920
rect 570328 26868 570380 26920
rect 145840 25712 145892 25764
rect 304356 25712 304408 25764
rect 151452 25644 151504 25696
rect 371700 25644 371752 25696
rect 160468 25576 160520 25628
rect 502984 25576 503036 25628
rect 20628 25508 20680 25560
rect 107016 25508 107068 25560
rect 161756 25508 161808 25560
rect 521844 25508 521896 25560
rect 140412 24420 140464 24472
rect 237012 24420 237064 24472
rect 147128 24352 147180 24404
rect 318524 24352 318576 24404
rect 152924 24284 152976 24336
rect 389456 24284 389508 24336
rect 168196 24216 168248 24268
rect 408408 24216 408460 24268
rect 160652 24148 160704 24200
rect 510068 24148 510120 24200
rect 163872 24080 163924 24132
rect 532516 24080 532568 24132
rect 144368 22856 144420 22908
rect 287796 22856 287848 22908
rect 168104 22788 168156 22840
rect 401324 22788 401376 22840
rect 161480 22720 161532 22772
rect 513564 22720 513616 22772
rect 140504 21632 140556 21684
rect 231032 21632 231084 21684
rect 148784 21564 148836 21616
rect 340972 21564 341024 21616
rect 148692 21496 148744 21548
rect 344560 21496 344612 21548
rect 149152 21428 149204 21480
rect 358728 21428 358780 21480
rect 133604 21360 133656 21412
rect 148324 21360 148376 21412
rect 149244 21360 149296 21412
rect 365812 21360 365864 21412
rect 143264 20204 143316 20256
rect 266544 20204 266596 20256
rect 144552 20136 144604 20188
rect 284300 20136 284352 20188
rect 144460 20068 144512 20120
rect 294880 20068 294932 20120
rect 159364 20000 159416 20052
rect 383568 20000 383620 20052
rect 169116 19932 169168 19984
rect 450912 19932 450964 19984
rect 137652 18776 137704 18828
rect 202696 18776 202748 18828
rect 139676 18708 139728 18760
rect 238116 18708 238168 18760
rect 151544 18640 151596 18692
rect 376484 18640 376536 18692
rect 11152 18572 11204 18624
rect 116860 18572 116912 18624
rect 166080 18572 166132 18624
rect 571524 18572 571576 18624
rect 138296 17484 138348 17536
rect 220452 17484 220504 17536
rect 168012 17416 168064 17468
rect 443828 17416 443880 17468
rect 157616 17348 157668 17400
rect 463976 17348 464028 17400
rect 157432 17280 157484 17332
rect 467472 17280 467524 17332
rect 43076 17212 43128 17264
rect 109684 17212 109736 17264
rect 132592 17212 132644 17264
rect 151084 17212 151136 17264
rect 157800 17212 157852 17264
rect 471060 17212 471112 17264
rect 138480 16124 138532 16176
rect 222752 16124 222804 16176
rect 147220 16056 147272 16108
rect 323308 16056 323360 16108
rect 150716 15988 150768 16040
rect 375288 15988 375340 16040
rect 150532 15920 150584 15972
rect 378876 15920 378928 15972
rect 35992 15852 36044 15904
rect 113916 15852 113968 15904
rect 152188 15852 152240 15904
rect 393044 15852 393096 15904
rect 143356 14696 143408 14748
rect 276020 14696 276072 14748
rect 144644 14628 144696 14680
rect 290188 14628 290240 14680
rect 148140 14560 148192 14612
rect 336280 14560 336332 14612
rect 167920 14492 167972 14544
rect 422576 14492 422628 14544
rect 28908 14424 28960 14476
rect 118148 14424 118200 14476
rect 154212 14424 154264 14476
rect 414296 14424 414348 14476
rect 139860 13336 139912 13388
rect 240508 13336 240560 13388
rect 147312 13268 147364 13320
rect 325608 13268 325660 13320
rect 154304 13200 154356 13252
rect 410800 13200 410852 13252
rect 155592 13132 155644 13184
rect 426164 13132 426216 13184
rect 85672 13064 85724 13116
rect 120908 13064 120960 13116
rect 133972 13064 134024 13116
rect 153844 13064 153896 13116
rect 165344 13064 165396 13116
rect 550272 13064 550324 13116
rect 132224 12384 132276 12436
rect 133144 12384 133196 12436
rect 167828 11772 167880 11824
rect 415492 11772 415544 11824
rect 158996 11704 159048 11756
rect 482836 11704 482888 11756
rect 147404 10480 147456 10532
rect 329196 10480 329248 10532
rect 155684 10412 155736 10464
rect 435548 10412 435600 10464
rect 46664 10344 46716 10396
rect 125508 10344 125560 10396
rect 169024 10344 169076 10396
rect 458088 10344 458140 10396
rect 19432 10276 19484 10328
rect 118056 10276 118108 10328
rect 163964 10276 164016 10328
rect 534908 10276 534960 10328
rect 145932 9256 145984 9308
rect 309048 9256 309100 9308
rect 145104 9188 145156 9240
rect 312636 9188 312688 9240
rect 149428 9120 149480 9172
rect 364616 9120 364668 9172
rect 154396 9052 154448 9104
rect 411904 9052 411956 9104
rect 159180 8984 159232 9036
rect 478144 8984 478196 9036
rect 96252 8916 96304 8968
rect 128912 8916 128964 8968
rect 164056 8916 164108 8968
rect 531320 8916 531372 8968
rect 471244 8236 471296 8288
rect 479340 8236 479392 8288
rect 142160 7760 142212 7812
rect 265348 7760 265400 7812
rect 147956 7692 148008 7744
rect 339868 7692 339920 7744
rect 50160 7624 50212 7676
rect 125416 7624 125468 7676
rect 155776 7624 155828 7676
rect 428464 7624 428516 7676
rect 24216 7556 24268 7608
rect 116768 7556 116820 7608
rect 163228 7556 163280 7608
rect 541992 7556 542044 7608
rect 141792 6808 141844 6860
rect 248788 6808 248840 6860
rect 141516 6740 141568 6792
rect 252376 6740 252428 6792
rect 141608 6672 141660 6724
rect 254676 6672 254728 6724
rect 141884 6604 141936 6656
rect 258264 6604 258316 6656
rect 141700 6536 141752 6588
rect 261760 6536 261812 6588
rect 2780 6468 2832 6520
rect 4804 6468 4856 6520
rect 145012 6468 145064 6520
rect 301964 6468 302016 6520
rect 145380 6400 145432 6452
rect 305552 6400 305604 6452
rect 153200 6332 153252 6384
rect 417884 6332 417936 6384
rect 154672 6264 154724 6316
rect 433248 6264 433300 6316
rect 78588 6196 78640 6248
rect 127440 6196 127492 6248
rect 132408 6196 132460 6248
rect 137652 6196 137704 6248
rect 164608 6196 164660 6248
rect 556160 6196 556212 6248
rect 6460 6128 6512 6180
rect 122196 6128 122248 6180
rect 122288 6128 122340 6180
rect 127624 6128 127676 6180
rect 132776 6128 132828 6180
rect 151820 6128 151872 6180
rect 164792 6128 164844 6180
rect 557356 6128 557408 6180
rect 136824 6060 136876 6112
rect 205088 6060 205140 6112
rect 137744 5992 137796 6044
rect 195612 5992 195664 6044
rect 132316 5516 132368 5568
rect 133788 5516 133840 5568
rect 137008 5108 137060 5160
rect 199108 5108 199160 5160
rect 146484 5040 146536 5092
rect 322112 5040 322164 5092
rect 147496 4972 147548 5024
rect 330392 4972 330444 5024
rect 157984 4904 158036 4956
rect 390652 4904 390704 4956
rect 71504 4836 71556 4888
rect 120724 4836 120776 4888
rect 152372 4836 152424 4888
rect 400128 4836 400180 4888
rect 5264 4768 5316 4820
rect 25504 4768 25556 4820
rect 45468 4768 45520 4820
rect 125232 4768 125284 4820
rect 134524 4768 134576 4820
rect 143540 4768 143592 4820
rect 166264 4768 166316 4820
rect 498200 4768 498252 4820
rect 141148 4088 141200 4140
rect 257068 4088 257120 4140
rect 141240 4020 141292 4072
rect 260656 4020 260708 4072
rect 151084 3952 151136 4004
rect 153016 3952 153068 4004
rect 160744 3952 160796 4004
rect 162492 3952 162544 4004
rect 167644 3952 167696 4004
rect 303160 3952 303212 4004
rect 144000 3884 144052 3936
rect 292580 3884 292632 3936
rect 108120 3816 108172 3868
rect 119344 3816 119396 3868
rect 170404 3816 170456 3868
rect 187332 3816 187384 3868
rect 189816 3816 189868 3868
rect 346952 3816 347004 3868
rect 98644 3748 98696 3800
rect 111064 3748 111116 3800
rect 136180 3748 136232 3800
rect 147128 3748 147180 3800
rect 156236 3748 156288 3800
rect 452108 3748 452160 3800
rect 66720 3680 66772 3732
rect 120816 3680 120868 3732
rect 134616 3680 134668 3732
rect 145932 3680 145984 3732
rect 167736 3680 167788 3732
rect 462780 3680 462832 3732
rect 51356 3612 51408 3664
rect 119528 3612 119580 3664
rect 135904 3612 135956 3664
rect 149520 3612 149572 3664
rect 151176 3612 151228 3664
rect 155408 3612 155460 3664
rect 156420 3612 156472 3664
rect 455696 3612 455748 3664
rect 475384 3612 475436 3664
rect 546684 3612 546736 3664
rect 15936 3544 15988 3596
rect 119436 3544 119488 3596
rect 135996 3544 136048 3596
rect 150624 3544 150676 3596
rect 156696 3544 156748 3596
rect 164884 3544 164936 3596
rect 173256 3544 173308 3596
rect 475752 3544 475804 3596
rect 508504 3544 508556 3596
rect 524236 3544 524288 3596
rect 1676 3476 1728 3528
rect 116676 3476 116728 3528
rect 125876 3476 125928 3528
rect 129004 3476 129056 3528
rect 129372 3476 129424 3528
rect 130660 3476 130712 3528
rect 134708 3476 134760 3528
rect 135260 3476 135312 3528
rect 136272 3476 136324 3528
rect 154212 3476 154264 3528
rect 155224 3476 155276 3528
rect 157800 3476 157852 3528
rect 162124 3476 162176 3528
rect 163688 3476 163740 3528
rect 170588 3476 170640 3528
rect 508872 3476 508924 3528
rect 572 3408 624 3460
rect 117964 3408 118016 3460
rect 119896 3408 119948 3460
rect 126244 3408 126296 3460
rect 126980 3408 127032 3460
rect 130476 3408 130528 3460
rect 130568 3408 130620 3460
rect 131948 3408 132000 3460
rect 133144 3408 133196 3460
rect 136456 3408 136508 3460
rect 17040 3340 17092 3392
rect 18604 3340 18656 3392
rect 37188 3340 37240 3392
rect 37924 3340 37976 3392
rect 69112 3340 69164 3392
rect 71044 3340 71096 3392
rect 110512 3340 110564 3392
rect 112444 3340 112496 3392
rect 134064 3340 134116 3392
rect 166080 3408 166132 3460
rect 170496 3408 170548 3460
rect 583392 3408 583444 3460
rect 184204 3340 184256 3392
rect 229836 3340 229888 3392
rect 153844 3272 153896 3324
rect 158904 3272 158956 3324
rect 577504 3272 577556 3324
rect 582196 3272 582248 3324
rect 104532 3204 104584 3256
rect 105544 3204 105596 3256
rect 111616 3204 111668 3256
rect 113824 3204 113876 3256
rect 39580 3068 39632 3120
rect 40776 3068 40828 3120
rect 178684 3068 178736 3120
rect 182548 3068 182600 3120
rect 27712 2932 27764 2984
rect 29644 2932 29696 2984
rect 124680 2932 124732 2984
rect 130384 2932 130436 2984
rect 136364 2932 136416 2984
rect 141240 2932 141292 2984
rect 158076 2932 158128 2984
rect 160100 2932 160152 2984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2778 449576 2834 449585
rect 2778 449511 2780 449520
rect 2832 449511 2834 449520
rect 2780 449482 2832 449488
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2792 345234 2820 345335
rect 2780 345228 2832 345234
rect 2780 345170 2832 345176
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3344 240174 3372 241023
rect 3332 240168 3384 240174
rect 3332 240110 3384 240116
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 210361 3372 214911
rect 3330 210352 3386 210361
rect 3330 210287 3386 210296
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3160 187746 3188 188799
rect 3148 187740 3200 187746
rect 3148 187682 3200 187688
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3344 162081 3372 162823
rect 3330 162072 3386 162081
rect 3330 162007 3386 162016
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3344 136678 3372 136711
rect 3332 136672 3384 136678
rect 3332 136614 3384 136620
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 3436 73137 3464 658135
rect 3698 566944 3754 566953
rect 3698 566879 3754 566888
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3422 73128 3478 73137
rect 3422 73063 3478 73072
rect 3528 70378 3556 501735
rect 3606 423600 3662 423609
rect 3606 423535 3662 423544
rect 3620 214849 3648 423535
rect 3712 384305 3740 566879
rect 4802 514856 4858 514865
rect 4802 514791 4858 514800
rect 3698 384296 3754 384305
rect 3698 384231 3754 384240
rect 3698 267200 3754 267209
rect 3698 267135 3754 267144
rect 3606 214840 3662 214849
rect 3606 214775 3662 214784
rect 3712 211857 3740 267135
rect 3698 211848 3754 211857
rect 3698 211783 3754 211792
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3620 133113 3648 149767
rect 3606 133104 3662 133113
rect 3606 133039 3662 133048
rect 3606 131200 3662 131209
rect 3606 131135 3662 131144
rect 3516 70372 3568 70378
rect 3516 70314 3568 70320
rect 2872 65544 2924 65550
rect 2872 65486 2924 65492
rect 2780 6520 2832 6526
rect 2778 6488 2780 6497
rect 2832 6488 2834 6497
rect 2778 6423 2834 6432
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 2884 480 2912 65486
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3422 33960 3478 33969
rect 3422 33895 3478 33904
rect 3436 32473 3464 33895
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3620 19417 3648 131135
rect 3698 128480 3754 128489
rect 3698 128415 3754 128424
rect 3712 58585 3740 128415
rect 3790 127120 3846 127129
rect 3790 127055 3846 127064
rect 3804 97617 3832 127055
rect 4816 117201 4844 514791
rect 4986 462632 5042 462641
rect 4986 462567 5042 462576
rect 4896 449540 4948 449546
rect 4896 449482 4948 449488
rect 4802 117192 4858 117201
rect 4802 117127 4858 117136
rect 3790 97608 3846 97617
rect 3790 97543 3846 97552
rect 4908 75546 4936 449482
rect 5000 118697 5028 462567
rect 5080 345228 5132 345234
rect 5080 345170 5132 345176
rect 4986 118688 5042 118697
rect 4986 118623 5042 118632
rect 4896 75540 4948 75546
rect 4896 75482 4948 75488
rect 5092 73778 5120 345170
rect 5080 73772 5132 73778
rect 5080 73714 5132 73720
rect 8128 73001 8156 703520
rect 15842 684312 15898 684321
rect 15842 684247 15898 684256
rect 11702 410544 11758 410553
rect 11702 410479 11758 410488
rect 11716 120057 11744 410479
rect 13084 397520 13136 397526
rect 13084 397462 13136 397468
rect 11702 120048 11758 120057
rect 11702 119983 11758 119992
rect 13096 75614 13124 397462
rect 14462 358456 14518 358465
rect 14462 358391 14518 358400
rect 14476 121417 14504 358391
rect 15856 136241 15884 684247
rect 18602 632088 18658 632097
rect 18602 632023 18658 632032
rect 18616 138689 18644 632023
rect 22742 580000 22798 580009
rect 22742 579935 22798 579944
rect 21364 240168 21416 240174
rect 21364 240110 21416 240116
rect 18602 138680 18658 138689
rect 18602 138615 18658 138624
rect 15842 136232 15898 136241
rect 15842 136167 15898 136176
rect 15842 134328 15898 134337
rect 15842 134263 15898 134272
rect 14462 121408 14518 121417
rect 14462 121343 14518 121352
rect 15856 110673 15884 134263
rect 17958 133104 18014 133113
rect 17958 133039 18014 133048
rect 17972 126993 18000 133039
rect 17958 126984 18014 126993
rect 17958 126919 18014 126928
rect 15842 110664 15898 110673
rect 15842 110599 15898 110608
rect 13084 75608 13136 75614
rect 13084 75550 13136 75556
rect 21376 74497 21404 240110
rect 22756 142905 22784 579935
rect 22834 254144 22890 254153
rect 22834 254079 22890 254088
rect 22742 142896 22798 142905
rect 22742 142831 22798 142840
rect 22848 124137 22876 254079
rect 22834 124128 22890 124137
rect 22834 124063 22890 124072
rect 24320 110401 24348 703520
rect 26882 671256 26938 671265
rect 26882 671191 26938 671200
rect 25502 475688 25558 475697
rect 25502 475623 25558 475632
rect 25516 145625 25544 475623
rect 25594 384296 25650 384305
rect 25594 384231 25650 384240
rect 25502 145616 25558 145625
rect 25502 145551 25558 145560
rect 25608 115841 25636 384231
rect 25594 115832 25650 115841
rect 25594 115767 25650 115776
rect 26896 111761 26924 671191
rect 29642 619168 29698 619177
rect 29642 619103 29698 619112
rect 26974 371376 27030 371385
rect 26974 371311 27030 371320
rect 26988 146985 27016 371311
rect 26974 146976 27030 146985
rect 26974 146911 27030 146920
rect 29656 113121 29684 619103
rect 31022 527912 31078 527921
rect 31022 527847 31078 527856
rect 29734 319288 29790 319297
rect 29734 319223 29790 319232
rect 29748 148345 29776 319223
rect 29734 148336 29790 148345
rect 29734 148271 29790 148280
rect 31036 144129 31064 527847
rect 31114 306232 31170 306241
rect 31114 306167 31170 306176
rect 31022 144120 31078 144129
rect 31022 144055 31078 144064
rect 31128 122777 31156 306167
rect 40512 141545 40540 703520
rect 45374 700632 45430 700641
rect 45374 700567 45430 700576
rect 44914 700496 44970 700505
rect 44914 700431 44970 700440
rect 43444 605872 43496 605878
rect 43444 605814 43496 605820
rect 40498 141536 40554 141545
rect 40498 141471 40554 141480
rect 31114 122768 31170 122777
rect 31114 122703 31170 122712
rect 29642 113112 29698 113121
rect 29642 113047 29698 113056
rect 26882 111752 26938 111761
rect 26882 111687 26938 111696
rect 24306 110392 24362 110401
rect 24306 110327 24362 110336
rect 21362 74488 21418 74497
rect 21362 74423 21418 74432
rect 8114 72992 8170 73001
rect 8114 72927 8170 72936
rect 43456 72865 43484 605814
rect 43536 553444 43588 553450
rect 43536 553386 43588 553392
rect 43442 72856 43498 72865
rect 43442 72791 43498 72800
rect 25502 72584 25558 72593
rect 25502 72519 25558 72528
rect 23020 72480 23072 72486
rect 23020 72422 23072 72428
rect 18234 71088 18290 71097
rect 18234 71023 18290 71032
rect 7656 68332 7708 68338
rect 7656 68274 7708 68280
rect 4804 63028 4856 63034
rect 4804 62970 4856 62976
rect 3698 58576 3754 58585
rect 3698 58511 3754 58520
rect 4068 46232 4120 46238
rect 4068 46174 4120 46180
rect 3606 19408 3662 19417
rect 3606 19343 3662 19352
rect 4080 480 4108 46174
rect 4816 6526 4844 62970
rect 4804 6520 4856 6526
rect 4804 6462 4856 6468
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5276 480 5304 4762
rect 6472 480 6500 6122
rect 7668 480 7696 68274
rect 12348 64184 12400 64190
rect 12348 64126 12400 64132
rect 9956 60036 10008 60042
rect 9956 59978 10008 59984
rect 8760 57248 8812 57254
rect 8760 57190 8812 57196
rect 8772 480 8800 57190
rect 9968 480 9996 59978
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 480 11192 18566
rect 12360 480 12388 64126
rect 13544 51740 13596 51746
rect 13544 51682 13596 51688
rect 13556 480 13584 51682
rect 14740 50380 14792 50386
rect 14740 50322 14792 50328
rect 14752 480 14780 50322
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15948 480 15976 3538
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 480 17080 3334
rect 18248 480 18276 71023
rect 21822 66872 21878 66881
rect 21822 66807 21878 66816
rect 18602 51776 18658 51785
rect 18602 51711 18658 51720
rect 18616 3398 18644 51711
rect 20628 25560 20680 25566
rect 20628 25502 20680 25508
rect 19432 10328 19484 10334
rect 19432 10270 19484 10276
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 19444 480 19472 10270
rect 20640 480 20668 25502
rect 21836 480 21864 66807
rect 23032 480 23060 72422
rect 25320 58676 25372 58682
rect 25320 58618 25372 58624
rect 24216 7608 24268 7614
rect 24216 7550 24268 7556
rect 24228 480 24256 7550
rect 25332 480 25360 58618
rect 25516 4826 25544 72519
rect 41880 71120 41932 71126
rect 41880 71062 41932 71068
rect 29644 71052 29696 71058
rect 29644 70994 29696 71000
rect 26516 65612 26568 65618
rect 26516 65554 26568 65560
rect 25504 4820 25556 4826
rect 25504 4762 25556 4768
rect 26528 480 26556 65554
rect 28908 14476 28960 14482
rect 28908 14418 28960 14424
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 27724 480 27752 2926
rect 28920 480 28948 14418
rect 29656 2990 29684 70994
rect 30104 68400 30156 68406
rect 30104 68342 30156 68348
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 30116 480 30144 68342
rect 34794 67008 34850 67017
rect 34794 66943 34850 66952
rect 32404 55888 32456 55894
rect 32404 55830 32456 55836
rect 31300 53100 31352 53106
rect 31300 53042 31352 53048
rect 31312 480 31340 53042
rect 32416 480 32444 55830
rect 33600 54528 33652 54534
rect 33600 54470 33652 54476
rect 33612 480 33640 54470
rect 34808 480 34836 66943
rect 40684 61396 40736 61402
rect 40684 61338 40736 61344
rect 38382 53136 38438 53145
rect 38382 53071 38438 53080
rect 37922 48920 37978 48929
rect 37922 48855 37978 48864
rect 35992 15904 36044 15910
rect 35992 15846 36044 15852
rect 36004 480 36032 15846
rect 37936 3398 37964 48855
rect 37188 3392 37240 3398
rect 37188 3334 37240 3340
rect 37924 3392 37976 3398
rect 37924 3334 37976 3340
rect 37200 480 37228 3334
rect 38396 480 38424 53071
rect 39580 3120 39632 3126
rect 39580 3062 39632 3068
rect 39592 480 39620 3062
rect 40696 480 40724 61338
rect 40774 50280 40830 50289
rect 40774 50215 40830 50224
rect 40788 3126 40816 50215
rect 40776 3120 40828 3126
rect 40776 3062 40828 3068
rect 41892 480 41920 71062
rect 43548 70310 43576 553386
rect 43628 292596 43680 292602
rect 43628 292538 43680 292544
rect 43640 75750 43668 292538
rect 44824 226024 44876 226030
rect 44824 225966 44876 225972
rect 44730 224224 44786 224233
rect 44730 224159 44786 224168
rect 44744 216209 44772 224159
rect 44730 216200 44786 216209
rect 44730 216135 44786 216144
rect 43628 75744 43680 75750
rect 43628 75686 43680 75692
rect 43536 70304 43588 70310
rect 44836 70281 44864 225966
rect 44928 106185 44956 700431
rect 45192 350124 45244 350130
rect 45192 350066 45244 350072
rect 45098 226128 45154 226137
rect 45098 226063 45154 226072
rect 45008 225004 45060 225010
rect 45008 224946 45060 224952
rect 45020 135930 45048 224946
rect 45008 135924 45060 135930
rect 45008 135866 45060 135872
rect 45112 109041 45140 226063
rect 45204 214606 45232 350066
rect 45284 249824 45336 249830
rect 45284 249766 45336 249772
rect 45296 215966 45324 249766
rect 45284 215960 45336 215966
rect 45284 215902 45336 215908
rect 45192 214600 45244 214606
rect 45192 214542 45244 214548
rect 45098 109032 45154 109041
rect 45098 108967 45154 108976
rect 45388 107545 45416 700567
rect 45742 700360 45798 700369
rect 45742 700295 45798 700304
rect 45468 224052 45520 224058
rect 45468 223994 45520 224000
rect 45480 209982 45508 223994
rect 45468 209976 45520 209982
rect 45468 209918 45520 209924
rect 45374 107536 45430 107545
rect 45374 107471 45430 107480
rect 44914 106176 44970 106185
rect 44914 106111 44970 106120
rect 45756 104825 45784 700295
rect 64144 413296 64196 413302
rect 64144 413238 64196 413244
rect 64156 405006 64184 413238
rect 50988 405000 51040 405006
rect 50988 404942 51040 404948
rect 64144 405000 64196 405006
rect 64144 404942 64196 404948
rect 51000 401674 51028 404942
rect 47584 401668 47636 401674
rect 47584 401610 47636 401616
rect 50988 401668 51040 401674
rect 50988 401610 51040 401616
rect 47596 382294 47624 401610
rect 46204 382288 46256 382294
rect 46204 382230 46256 382236
rect 47584 382288 47636 382294
rect 47584 382230 47636 382236
rect 46216 350130 46244 382230
rect 58624 356720 58676 356726
rect 58624 356662 58676 356668
rect 46204 350124 46256 350130
rect 46204 350066 46256 350072
rect 58636 339726 58664 356662
rect 57244 339720 57296 339726
rect 57244 339662 57296 339668
rect 58624 339720 58676 339726
rect 58624 339662 58676 339668
rect 57256 327078 57284 339662
rect 55956 327072 56008 327078
rect 55956 327014 56008 327020
rect 57244 327072 57296 327078
rect 57244 327014 57296 327020
rect 55968 321162 55996 327014
rect 54484 321156 54536 321162
rect 54484 321098 54536 321104
rect 55956 321156 56008 321162
rect 55956 321098 56008 321104
rect 54496 309126 54524 321098
rect 53104 309120 53156 309126
rect 53104 309062 53156 309068
rect 54484 309120 54536 309126
rect 54484 309062 54536 309068
rect 53116 279478 53144 309062
rect 70950 281616 71006 281625
rect 70950 281551 71006 281560
rect 57888 280832 57940 280838
rect 57888 280774 57940 280780
rect 51080 279472 51132 279478
rect 51080 279414 51132 279420
rect 53104 279472 53156 279478
rect 53104 279414 53156 279420
rect 47584 278044 47636 278050
rect 47584 277986 47636 277992
rect 47596 270230 47624 277986
rect 51092 277394 51120 279414
rect 57900 278050 57928 280774
rect 70964 280129 70992 281551
rect 69662 280120 69718 280129
rect 69662 280055 69718 280064
rect 70950 280120 71006 280129
rect 70950 280055 71006 280064
rect 57888 278044 57940 278050
rect 57888 277986 57940 277992
rect 51000 277366 51120 277394
rect 51000 273290 51028 277366
rect 69676 276049 69704 280055
rect 67822 276040 67878 276049
rect 67822 275975 67878 275984
rect 69662 276040 69718 276049
rect 69662 275975 69718 275984
rect 48964 273284 49016 273290
rect 48964 273226 49016 273232
rect 50988 273284 51040 273290
rect 50988 273226 51040 273232
rect 46204 270224 46256 270230
rect 46204 270166 46256 270172
rect 47584 270224 47636 270230
rect 47584 270166 47636 270172
rect 45834 224904 45890 224913
rect 45834 224839 45890 224848
rect 45848 215937 45876 224839
rect 46216 224058 46244 270166
rect 48976 262274 49004 273226
rect 67836 270473 67864 275975
rect 66534 270464 66590 270473
rect 66534 270399 66590 270408
rect 67822 270464 67878 270473
rect 67822 270399 67878 270408
rect 66548 265033 66576 270399
rect 65522 265024 65578 265033
rect 65522 264959 65578 264968
rect 66534 265024 66590 265033
rect 66534 264959 66590 264968
rect 47676 262268 47728 262274
rect 47676 262210 47728 262216
rect 48964 262268 49016 262274
rect 48964 262210 49016 262216
rect 47688 259282 47716 262210
rect 46296 259276 46348 259282
rect 46296 259218 46348 259224
rect 47676 259276 47728 259282
rect 47676 259218 47728 259224
rect 46308 249830 46336 259218
rect 46296 249824 46348 249830
rect 46296 249766 46348 249772
rect 65536 248441 65564 264959
rect 64142 248432 64198 248441
rect 64142 248367 64198 248376
rect 65522 248432 65578 248441
rect 65522 248367 65578 248376
rect 64156 231169 64184 248367
rect 53838 231160 53894 231169
rect 53838 231095 53894 231104
rect 64142 231160 64198 231169
rect 64142 231095 64198 231104
rect 53852 225049 53880 231095
rect 68926 226264 68982 226273
rect 68926 226199 68982 226208
rect 53838 225040 53894 225049
rect 68940 225010 68968 226199
rect 72988 226030 73016 703520
rect 79324 436756 79376 436762
rect 79324 436698 79376 436704
rect 79336 419558 79364 436698
rect 76932 419552 76984 419558
rect 76932 419494 76984 419500
rect 79324 419552 79376 419558
rect 79324 419494 79376 419500
rect 76944 417858 76972 419494
rect 73160 417852 73212 417858
rect 73160 417794 73212 417800
rect 76932 417852 76984 417858
rect 76932 417794 76984 417800
rect 73172 413302 73200 417794
rect 73160 413296 73212 413302
rect 73160 413238 73212 413244
rect 77942 334656 77998 334665
rect 77942 334591 77998 334600
rect 77956 320929 77984 334591
rect 76562 320920 76618 320929
rect 76562 320855 76618 320864
rect 77942 320920 77998 320929
rect 77942 320855 77998 320864
rect 76576 291145 76604 320855
rect 87604 305040 87656 305046
rect 87604 304982 87656 304988
rect 75274 291136 75330 291145
rect 75274 291071 75330 291080
rect 76562 291136 76618 291145
rect 76562 291071 76618 291080
rect 75288 288561 75316 291071
rect 73250 288552 73306 288561
rect 73250 288487 73306 288496
rect 75274 288552 75330 288561
rect 75274 288487 75330 288496
rect 73160 287700 73212 287706
rect 73160 287642 73212 287648
rect 73172 280838 73200 287642
rect 73264 281625 73292 288487
rect 87616 287706 87644 304982
rect 87604 287700 87656 287706
rect 87604 287642 87656 287648
rect 73250 281616 73306 281625
rect 73250 281551 73306 281560
rect 73160 280832 73212 280838
rect 73160 280774 73212 280780
rect 89180 226137 89208 703520
rect 93124 461644 93176 461650
rect 93124 461586 93176 461592
rect 93136 436762 93164 461586
rect 93124 436756 93176 436762
rect 93124 436698 93176 436704
rect 95240 337408 95292 337414
rect 95240 337350 95292 337356
rect 95252 328914 95280 337350
rect 93124 328908 93176 328914
rect 93124 328850 93176 328856
rect 95240 328908 95292 328914
rect 95240 328850 95292 328856
rect 93136 305046 93164 328850
rect 93124 305040 93176 305046
rect 93124 304982 93176 304988
rect 98918 236736 98974 236745
rect 98918 236671 98974 236680
rect 98932 230489 98960 236671
rect 95238 230480 95294 230489
rect 95238 230415 95294 230424
rect 98918 230480 98974 230489
rect 98918 230415 98974 230424
rect 89166 226128 89222 226137
rect 89166 226063 89222 226072
rect 72976 226024 73028 226030
rect 72976 225966 73028 225972
rect 53838 224975 53894 224984
rect 68928 225004 68980 225010
rect 68928 224946 68980 224952
rect 95252 224233 95280 230415
rect 105464 226273 105492 703520
rect 134800 574116 134852 574122
rect 134800 574058 134852 574064
rect 134812 570994 134840 574058
rect 127624 570988 127676 570994
rect 127624 570930 127676 570936
rect 134800 570988 134852 570994
rect 134800 570930 134852 570936
rect 127636 552702 127664 570930
rect 124864 552696 124916 552702
rect 124864 552638 124916 552644
rect 127624 552696 127676 552702
rect 127624 552638 127676 552644
rect 124876 532098 124904 552638
rect 119344 532092 119396 532098
rect 119344 532034 119396 532040
rect 124864 532092 124916 532098
rect 124864 532034 124916 532040
rect 119356 511222 119384 532034
rect 114560 511216 114612 511222
rect 114560 511158 114612 511164
rect 119344 511216 119396 511222
rect 119344 511158 119396 511164
rect 114572 504218 114600 511158
rect 137848 508570 137876 703520
rect 154132 700641 154160 703520
rect 154118 700632 154174 700641
rect 154118 700567 154174 700576
rect 156604 643748 156656 643754
rect 156604 643690 156656 643696
rect 156616 635526 156644 643690
rect 150440 635520 150492 635526
rect 150440 635462 150492 635468
rect 156604 635520 156656 635526
rect 156604 635462 156656 635468
rect 150452 631378 150480 635462
rect 141424 631372 141476 631378
rect 141424 631314 141476 631320
rect 150440 631372 150492 631378
rect 150440 631314 150492 631320
rect 141436 574122 141464 631314
rect 141424 574116 141476 574122
rect 141424 574058 141476 574064
rect 117964 508564 118016 508570
rect 117964 508506 118016 508512
rect 137836 508564 137888 508570
rect 137836 508506 137888 508512
rect 112444 504212 112496 504218
rect 112444 504154 112496 504160
rect 114560 504212 114612 504218
rect 114560 504154 114612 504160
rect 112456 461650 112484 504154
rect 117976 487218 118004 508506
rect 116584 487212 116636 487218
rect 116584 487154 116636 487160
rect 117964 487212 118016 487218
rect 117964 487154 118016 487160
rect 116596 473006 116624 487154
rect 115204 473000 115256 473006
rect 115204 472942 115256 472948
rect 116584 473000 116636 473006
rect 116584 472942 116636 472948
rect 112444 461644 112496 461650
rect 112444 461586 112496 461592
rect 115216 356726 115244 472942
rect 166264 467152 166316 467158
rect 166264 467094 166316 467100
rect 166276 452878 166304 467094
rect 162860 452872 162912 452878
rect 162860 452814 162912 452820
rect 166264 452872 166316 452878
rect 166264 452814 166316 452820
rect 162872 447098 162900 452814
rect 155224 447092 155276 447098
rect 155224 447034 155276 447040
rect 162860 447092 162912 447098
rect 162860 447034 162912 447040
rect 155236 411330 155264 447034
rect 167642 440872 167698 440881
rect 167642 440807 167698 440816
rect 167656 427961 167684 440807
rect 164882 427952 164938 427961
rect 164882 427887 164938 427896
rect 167642 427952 167698 427961
rect 167642 427887 167698 427896
rect 152464 411324 152516 411330
rect 152464 411266 152516 411272
rect 155224 411324 155276 411330
rect 155224 411266 155276 411272
rect 152476 363662 152504 411266
rect 115296 363656 115348 363662
rect 115296 363598 115348 363604
rect 152464 363656 152516 363662
rect 152464 363598 152516 363604
rect 115204 356720 115256 356726
rect 115204 356662 115256 356668
rect 115308 337414 115336 363598
rect 164896 356697 164924 427887
rect 153842 356688 153898 356697
rect 153842 356623 153898 356632
rect 164882 356688 164938 356697
rect 164882 356623 164938 356632
rect 153856 342145 153884 356623
rect 145838 342136 145894 342145
rect 145838 342071 145894 342080
rect 153842 342136 153898 342145
rect 153842 342071 153898 342080
rect 145852 338065 145880 342071
rect 142802 338056 142858 338065
rect 142802 337991 142858 338000
rect 145838 338056 145894 338065
rect 145838 337991 145894 338000
rect 115296 337408 115348 337414
rect 115296 337350 115348 337356
rect 142816 323649 142844 337991
rect 170324 334665 170352 703520
rect 202800 700058 202828 703520
rect 218992 700505 219020 703520
rect 235184 700505 235212 703520
rect 218978 700496 219034 700505
rect 218978 700431 219034 700440
rect 220082 700496 220138 700505
rect 220082 700431 220138 700440
rect 235170 700496 235226 700505
rect 235170 700431 235226 700440
rect 194692 700052 194744 700058
rect 194692 699994 194744 700000
rect 202788 700052 202840 700058
rect 202788 699994 202840 700000
rect 194704 696998 194732 699994
rect 193128 696992 193180 696998
rect 193128 696934 193180 696940
rect 194692 696992 194744 696998
rect 194692 696934 194744 696940
rect 193140 694210 193168 696934
rect 188344 694204 188396 694210
rect 188344 694146 188396 694152
rect 193128 694204 193180 694210
rect 193128 694146 193180 694152
rect 188356 679114 188384 694146
rect 183192 679108 183244 679114
rect 183192 679050 183244 679056
rect 188344 679108 188396 679114
rect 188344 679050 188396 679056
rect 183204 677210 183232 679050
rect 180064 677204 180116 677210
rect 180064 677146 180116 677152
rect 183192 677204 183244 677210
rect 183192 677146 183244 677152
rect 180076 657218 180104 677146
rect 175924 657212 175976 657218
rect 175924 657154 175976 657160
rect 180064 657212 180116 657218
rect 180064 657154 180116 657160
rect 175936 643754 175964 657154
rect 220096 644609 220124 700431
rect 267660 699718 267688 703520
rect 283852 700369 283880 703520
rect 283838 700360 283894 700369
rect 283838 700295 283894 700304
rect 300136 699961 300164 703520
rect 332520 700330 332548 703520
rect 348804 700369 348832 703520
rect 364996 700505 365024 703520
rect 364982 700496 365038 700505
rect 364982 700431 365038 700440
rect 396538 700496 396594 700505
rect 396538 700431 396594 700440
rect 348790 700360 348846 700369
rect 332508 700324 332560 700330
rect 348790 700295 348846 700304
rect 332508 700266 332560 700272
rect 300122 699952 300178 699961
rect 300122 699887 300178 699896
rect 303158 699952 303214 699961
rect 303158 699887 303214 699896
rect 260104 699712 260156 699718
rect 260104 699654 260156 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 260116 690334 260144 699654
rect 303172 697513 303200 699887
rect 303158 697504 303214 697513
rect 303158 697439 303214 697448
rect 309782 697504 309838 697513
rect 309782 697439 309838 697448
rect 253940 690328 253992 690334
rect 253940 690270 253992 690276
rect 260104 690328 260156 690334
rect 260104 690270 260156 690276
rect 253952 683806 253980 690270
rect 309796 690169 309824 697439
rect 309782 690160 309838 690169
rect 309782 690095 309838 690104
rect 312542 690160 312598 690169
rect 312542 690095 312598 690104
rect 312556 685817 312584 690095
rect 312542 685808 312598 685817
rect 312542 685743 312598 685752
rect 315302 685808 315358 685817
rect 315302 685743 315358 685752
rect 238760 683800 238812 683806
rect 238760 683742 238812 683748
rect 253940 683800 253992 683806
rect 253940 683742 253992 683748
rect 238772 679930 238800 683742
rect 233884 679924 233936 679930
rect 233884 679866 233936 679872
rect 238760 679924 238812 679930
rect 238760 679866 238812 679872
rect 213182 644600 213238 644609
rect 213182 644535 213238 644544
rect 220082 644600 220138 644609
rect 220082 644535 220138 644544
rect 175924 643748 175976 643754
rect 175924 643690 175976 643696
rect 211804 591320 211856 591326
rect 211804 591262 211856 591268
rect 207662 589928 207718 589937
rect 207662 589863 207718 589872
rect 195244 570648 195296 570654
rect 195244 570590 195296 570596
rect 195256 567866 195284 570590
rect 189724 567860 189776 567866
rect 189724 567802 189776 567808
rect 195244 567860 195296 567866
rect 195244 567802 195296 567808
rect 189736 511970 189764 567802
rect 207676 551993 207704 589863
rect 211816 580990 211844 591262
rect 213196 589937 213224 644535
rect 233896 591326 233924 679866
rect 315316 663921 315344 685743
rect 315302 663912 315358 663921
rect 315302 663847 315358 663856
rect 317418 663912 317474 663921
rect 317418 663847 317474 663856
rect 317432 658889 317460 663847
rect 317418 658880 317474 658889
rect 317418 658815 317474 658824
rect 337382 658880 337438 658889
rect 337382 658815 337438 658824
rect 337396 646513 337424 658815
rect 337382 646504 337438 646513
rect 337382 646439 337438 646448
rect 345018 646504 345074 646513
rect 345018 646439 345074 646448
rect 345032 639713 345060 646439
rect 345018 639704 345074 639713
rect 345018 639639 345074 639648
rect 348422 639704 348478 639713
rect 348422 639639 348478 639648
rect 233884 591320 233936 591326
rect 233884 591262 233936 591268
rect 213182 589928 213238 589937
rect 213182 589863 213238 589872
rect 209044 580984 209096 580990
rect 209044 580926 209096 580932
rect 211804 580984 211856 580990
rect 211804 580926 211856 580932
rect 209056 570654 209084 580926
rect 209044 570648 209096 570654
rect 209044 570590 209096 570596
rect 204902 551984 204958 551993
rect 204902 551919 204958 551928
rect 207662 551984 207718 551993
rect 207662 551919 207718 551928
rect 184388 511964 184440 511970
rect 184388 511906 184440 511912
rect 189724 511964 189776 511970
rect 189724 511906 189776 511912
rect 184400 507142 184428 511906
rect 178684 507136 178736 507142
rect 178684 507078 178736 507084
rect 184388 507136 184440 507142
rect 184388 507078 184440 507084
rect 178696 483002 178724 507078
rect 174544 482996 174596 483002
rect 174544 482938 174596 482944
rect 178684 482996 178736 483002
rect 178684 482938 178736 482944
rect 174556 467158 174584 482938
rect 204916 480865 204944 551919
rect 348436 525881 348464 639639
rect 348422 525872 348478 525881
rect 348422 525807 348478 525816
rect 351182 525872 351238 525881
rect 351182 525807 351238 525816
rect 197266 480856 197322 480865
rect 197266 480791 197322 480800
rect 204902 480856 204958 480865
rect 204902 480791 204958 480800
rect 197280 478145 197308 480791
rect 184202 478136 184258 478145
rect 184202 478071 184258 478080
rect 197266 478136 197322 478145
rect 197266 478071 197322 478080
rect 174544 467152 174596 467158
rect 174544 467094 174596 467100
rect 184216 457473 184244 478071
rect 178682 457464 178738 457473
rect 178682 457399 178738 457408
rect 184202 457464 184258 457473
rect 184202 457399 184258 457408
rect 178696 440881 178724 457399
rect 178682 440872 178738 440881
rect 178682 440807 178738 440816
rect 351196 351121 351224 525807
rect 351182 351112 351238 351121
rect 351182 351047 351238 351056
rect 376022 351112 376078 351121
rect 376022 351047 376078 351056
rect 376036 339425 376064 351047
rect 376022 339416 376078 339425
rect 376022 339351 376078 339360
rect 378782 339416 378838 339425
rect 378782 339351 378838 339360
rect 170310 334656 170366 334665
rect 170310 334591 170366 334600
rect 378796 332489 378824 339351
rect 378782 332480 378838 332489
rect 378782 332415 378838 332424
rect 384578 332480 384634 332489
rect 384578 332415 384634 332424
rect 384592 329089 384620 332415
rect 384578 329080 384634 329089
rect 384578 329015 384634 329024
rect 395342 329080 395398 329089
rect 395342 329015 395398 329024
rect 139398 323640 139454 323649
rect 139398 323575 139454 323584
rect 142802 323640 142858 323649
rect 142802 323575 142858 323584
rect 139412 316713 139440 323575
rect 129002 316704 129058 316713
rect 129002 316639 129058 316648
rect 139398 316704 139454 316713
rect 139398 316639 139454 316648
rect 129016 301617 129044 316639
rect 126242 301608 126298 301617
rect 126242 301543 126298 301552
rect 129002 301608 129058 301617
rect 129002 301543 129058 301552
rect 126256 287745 126284 301543
rect 120814 287736 120870 287745
rect 120814 287671 120870 287680
rect 126242 287736 126298 287745
rect 126242 287671 126298 287680
rect 120828 282305 120856 287671
rect 395356 285705 395384 329015
rect 395342 285696 395398 285705
rect 395342 285631 395398 285640
rect 396446 285696 396502 285705
rect 396446 285631 396502 285640
rect 117962 282296 118018 282305
rect 117962 282231 118018 282240
rect 120814 282296 120870 282305
rect 120814 282231 120870 282240
rect 117976 272241 118004 282231
rect 113822 272232 113878 272241
rect 113822 272167 113878 272176
rect 117962 272232 118018 272241
rect 117962 272167 118018 272176
rect 113836 266393 113864 272167
rect 108302 266384 108358 266393
rect 108302 266319 108358 266328
rect 113822 266384 113878 266393
rect 113822 266319 113878 266328
rect 108316 254017 108344 266319
rect 105542 254008 105598 254017
rect 105542 253943 105598 253952
rect 108302 254008 108358 254017
rect 108302 253943 108358 253952
rect 105556 236745 105584 253943
rect 105542 236736 105598 236745
rect 105542 236671 105598 236680
rect 105450 226264 105506 226273
rect 105450 226199 105506 226208
rect 95238 224224 95294 224233
rect 95238 224159 95294 224168
rect 46204 224052 46256 224058
rect 46204 223994 46256 224000
rect 46846 216200 46902 216209
rect 46846 216135 46902 216144
rect 45834 215928 45890 215937
rect 45834 215863 45890 215872
rect 46860 210497 46888 216135
rect 56692 215960 56744 215966
rect 57336 215960 57388 215966
rect 56744 215908 57336 215914
rect 56692 215902 57388 215908
rect 68284 215960 68336 215966
rect 68284 215902 68336 215908
rect 149058 215928 149114 215937
rect 56704 215886 57376 215902
rect 57730 214526 57928 214554
rect 57796 214328 57848 214334
rect 57796 214270 57848 214276
rect 46846 210488 46902 210497
rect 46846 210423 46902 210432
rect 56598 210488 56654 210497
rect 56598 210423 56654 210432
rect 47584 209976 47636 209982
rect 47584 209918 47636 209924
rect 47596 202842 47624 209918
rect 56612 205737 56640 210423
rect 57808 209098 57836 214270
rect 57796 209092 57848 209098
rect 57796 209034 57848 209040
rect 56598 205728 56654 205737
rect 56598 205663 56654 205672
rect 47584 202836 47636 202842
rect 47584 202778 47636 202784
rect 51724 202836 51776 202842
rect 51724 202778 51776 202784
rect 46202 201920 46258 201929
rect 46202 201855 46258 201864
rect 46216 125497 46244 201855
rect 51736 164898 51764 202778
rect 57900 193905 57928 214526
rect 68296 208962 68324 215902
rect 149058 215863 149114 215872
rect 114374 214704 114430 214713
rect 114374 214639 114430 214648
rect 87722 214526 88288 214554
rect 69664 209092 69716 209098
rect 69664 209034 69716 209040
rect 68284 208956 68336 208962
rect 68284 208898 68336 208904
rect 58622 205728 58678 205737
rect 58622 205663 58678 205672
rect 57886 193896 57942 193905
rect 57886 193831 57942 193840
rect 58636 191729 58664 205663
rect 69676 204950 69704 209034
rect 75552 208956 75604 208962
rect 75552 208898 75604 208904
rect 69664 204944 69716 204950
rect 69664 204886 69716 204892
rect 75564 201550 75592 208898
rect 85120 204944 85172 204950
rect 85120 204886 85172 204892
rect 75552 201544 75604 201550
rect 75552 201486 75604 201492
rect 85132 201482 85160 204886
rect 78036 201476 78088 201482
rect 78036 201418 78088 201424
rect 85120 201476 85172 201482
rect 85120 201418 85172 201424
rect 87604 201476 87656 201482
rect 87604 201418 87656 201424
rect 78048 198762 78076 201418
rect 78036 198756 78088 198762
rect 78036 198698 78088 198704
rect 81440 198688 81492 198694
rect 81440 198630 81492 198636
rect 81452 194614 81480 198630
rect 81440 194608 81492 194614
rect 81440 194550 81492 194556
rect 87616 194546 87644 201418
rect 84844 194540 84896 194546
rect 84844 194482 84896 194488
rect 87604 194540 87656 194546
rect 87604 194482 87656 194488
rect 58622 191720 58678 191729
rect 58622 191655 58678 191664
rect 60002 191720 60058 191729
rect 60002 191655 60058 191664
rect 60016 186425 60044 191655
rect 60002 186416 60058 186425
rect 60002 186351 60058 186360
rect 61382 186416 61438 186425
rect 61382 186351 61438 186360
rect 61396 167113 61424 186351
rect 84856 184890 84884 194482
rect 84844 184884 84896 184890
rect 84844 184826 84896 184832
rect 86224 184884 86276 184890
rect 86224 184826 86276 184832
rect 86236 179450 86264 184826
rect 88260 182073 88288 214526
rect 89720 194540 89772 194546
rect 89720 194482 89772 194488
rect 89732 191146 89760 194482
rect 89720 191140 89772 191146
rect 89720 191082 89772 191088
rect 111064 191140 111116 191146
rect 111064 191082 111116 191088
rect 111076 182782 111104 191082
rect 112444 187740 112496 187746
rect 112444 187682 112496 187688
rect 111064 182776 111116 182782
rect 111064 182718 111116 182724
rect 88246 182064 88302 182073
rect 88246 181999 88302 182008
rect 86224 179444 86276 179450
rect 86224 179386 86276 179392
rect 89444 179376 89496 179382
rect 89444 179318 89496 179324
rect 89456 173874 89484 179318
rect 89444 173868 89496 173874
rect 89444 173810 89496 173816
rect 92480 173868 92532 173874
rect 92480 173810 92532 173816
rect 61382 167104 61438 167113
rect 61382 167039 61438 167048
rect 62762 167104 62818 167113
rect 92492 167074 92520 173810
rect 62762 167039 62818 167048
rect 92480 167068 92532 167074
rect 51724 164892 51776 164898
rect 51724 164834 51776 164840
rect 62776 144265 62804 167039
rect 92480 167010 92532 167016
rect 95884 167000 95936 167006
rect 95884 166942 95936 166948
rect 66904 164892 66956 164898
rect 66904 164834 66956 164840
rect 66916 155922 66944 164834
rect 95896 155922 95924 166942
rect 66904 155916 66956 155922
rect 66904 155858 66956 155864
rect 69296 155916 69348 155922
rect 69296 155858 69348 155864
rect 95884 155916 95936 155922
rect 95884 155858 95936 155864
rect 97264 155916 97316 155922
rect 97264 155858 97316 155864
rect 69308 152522 69336 155858
rect 69296 152516 69348 152522
rect 69296 152458 69348 152464
rect 84200 152516 84252 152522
rect 84200 152458 84252 152464
rect 84212 149122 84240 152458
rect 84200 149116 84252 149122
rect 84200 149058 84252 149064
rect 87604 149116 87656 149122
rect 87604 149058 87656 149064
rect 62762 144256 62818 144265
rect 62762 144191 62818 144200
rect 70766 144256 70822 144265
rect 70766 144191 70822 144200
rect 70780 140865 70808 144191
rect 70766 140856 70822 140865
rect 70766 140791 70822 140800
rect 73158 140856 73214 140865
rect 73158 140791 73214 140800
rect 73172 134473 73200 140791
rect 73158 134464 73214 134473
rect 73158 134399 73214 134408
rect 46202 125488 46258 125497
rect 46202 125423 46258 125432
rect 87616 104854 87644 149058
rect 97276 129130 97304 155858
rect 97264 129124 97316 129130
rect 97264 129066 97316 129072
rect 102784 129124 102836 129130
rect 102784 129066 102836 129072
rect 102796 117366 102824 129066
rect 102784 117360 102836 117366
rect 102784 117302 102836 117308
rect 105544 117292 105596 117298
rect 105544 117234 105596 117240
rect 87604 104848 87656 104854
rect 45742 104816 45798 104825
rect 87604 104790 87656 104796
rect 90364 104848 90416 104854
rect 90364 104790 90416 104796
rect 45742 104751 45798 104760
rect 90376 100026 90404 104790
rect 90364 100020 90416 100026
rect 90364 99962 90416 99968
rect 101404 100020 101456 100026
rect 101404 99962 101456 99968
rect 101416 89690 101444 99962
rect 105556 92546 105584 117234
rect 105544 92540 105596 92546
rect 105544 92482 105596 92488
rect 109408 92540 109460 92546
rect 109408 92482 109460 92488
rect 109420 89758 109448 92482
rect 109408 89752 109460 89758
rect 109408 89694 109460 89700
rect 101404 89684 101456 89690
rect 101404 89626 101456 89632
rect 104164 89684 104216 89690
rect 104164 89626 104216 89632
rect 84476 71188 84528 71194
rect 84476 71130 84528 71136
rect 43536 70246 43588 70252
rect 44822 70272 44878 70281
rect 44822 70207 44878 70216
rect 80888 69896 80940 69902
rect 80888 69838 80940 69844
rect 71044 69828 71096 69834
rect 71044 69770 71096 69776
rect 54944 69760 54996 69766
rect 54944 69702 54996 69708
rect 47860 69692 47912 69698
rect 47860 69634 47912 69640
rect 44272 62824 44324 62830
rect 44272 62766 44324 62772
rect 43076 17264 43128 17270
rect 43076 17206 43128 17212
rect 43088 480 43116 17206
rect 44284 480 44312 62766
rect 46664 10396 46716 10402
rect 46664 10338 46716 10344
rect 45468 4820 45520 4826
rect 45468 4762 45520 4768
rect 45480 480 45508 4762
rect 46676 480 46704 10338
rect 47872 480 47900 69634
rect 48964 64252 49016 64258
rect 48964 64194 49016 64200
rect 48976 480 49004 64194
rect 52550 64152 52606 64161
rect 52550 64087 52606 64096
rect 50160 7676 50212 7682
rect 50160 7618 50212 7624
rect 50172 480 50200 7618
rect 51356 3664 51408 3670
rect 51356 3606 51408 3612
rect 51368 480 51396 3606
rect 52564 480 52592 64087
rect 53746 46200 53802 46209
rect 53746 46135 53802 46144
rect 53760 480 53788 46135
rect 54956 480 54984 69702
rect 58440 68468 58492 68474
rect 58440 68410 58492 68416
rect 56048 62892 56100 62898
rect 56048 62834 56100 62840
rect 56060 480 56088 62834
rect 57244 55956 57296 55962
rect 57244 55898 57296 55904
rect 57256 480 57284 55898
rect 58452 480 58480 68410
rect 60832 66904 60884 66910
rect 60832 66846 60884 66852
rect 59636 60104 59688 60110
rect 59636 60046 59688 60052
rect 59648 480 59676 60046
rect 60844 480 60872 66846
rect 67916 64320 67968 64326
rect 67916 64262 67968 64268
rect 65524 61464 65576 61470
rect 65524 61406 65576 61412
rect 63224 60172 63276 60178
rect 63224 60114 63276 60120
rect 62028 53168 62080 53174
rect 62028 53110 62080 53116
rect 62040 480 62068 53110
rect 63236 480 63264 60114
rect 64328 44872 64380 44878
rect 64328 44814 64380 44820
rect 64340 480 64368 44814
rect 65536 480 65564 61406
rect 66720 3732 66772 3738
rect 66720 3674 66772 3680
rect 66732 480 66760 3674
rect 67928 480 67956 64262
rect 70306 58712 70362 58721
rect 70306 58647 70362 58656
rect 69112 3392 69164 3398
rect 69112 3334 69164 3340
rect 69124 480 69152 3334
rect 70320 480 70348 58647
rect 71056 3398 71084 69770
rect 72606 68232 72662 68241
rect 72606 68167 72662 68176
rect 71504 4888 71556 4894
rect 71504 4830 71556 4836
rect 71044 3392 71096 3398
rect 71044 3334 71096 3340
rect 71516 480 71544 4830
rect 72620 480 72648 68167
rect 76196 66972 76248 66978
rect 76196 66914 76248 66920
rect 73802 50416 73858 50425
rect 73802 50351 73858 50360
rect 73816 480 73844 50351
rect 74998 49056 75054 49065
rect 74998 48991 75054 49000
rect 75012 480 75040 48991
rect 76208 480 76236 66914
rect 79692 65680 79744 65686
rect 79692 65622 79744 65628
rect 77392 57316 77444 57322
rect 77392 57258 77444 57264
rect 77404 480 77432 57258
rect 78588 6248 78640 6254
rect 78588 6190 78640 6196
rect 78600 480 78628 6190
rect 79704 480 79732 65622
rect 80900 480 80928 69838
rect 83280 47592 83332 47598
rect 83280 47534 83332 47540
rect 82084 40724 82136 40730
rect 82084 40666 82136 40672
rect 82096 480 82124 40666
rect 83292 480 83320 47534
rect 84488 480 84516 71130
rect 104176 70145 104204 89626
rect 112456 74254 112484 187682
rect 113548 182776 113600 182782
rect 113548 182718 113600 182724
rect 113560 180742 113588 182718
rect 113824 181144 113876 181150
rect 113824 181086 113876 181092
rect 113548 180736 113600 180742
rect 113548 180678 113600 180684
rect 113730 137320 113786 137329
rect 113730 137255 113786 137264
rect 112536 136672 112588 136678
rect 112536 136614 112588 136620
rect 112548 74390 112576 136614
rect 113744 91089 113772 137255
rect 113836 133249 113864 181086
rect 114006 156632 114062 156641
rect 114006 156567 114062 156576
rect 113914 142760 113970 142769
rect 113914 142695 113970 142704
rect 113822 133240 113878 133249
rect 113822 133175 113878 133184
rect 113822 129840 113878 129849
rect 113822 129775 113878 129784
rect 113730 91080 113786 91089
rect 113730 91015 113786 91024
rect 113836 80889 113864 129775
rect 113928 89729 113956 142695
rect 113914 89720 113970 89729
rect 113914 89655 113970 89664
rect 114020 88233 114048 156567
rect 114098 155272 114154 155281
rect 114098 155207 114154 155216
rect 114006 88224 114062 88233
rect 114006 88159 114062 88168
rect 114112 86873 114140 155207
rect 114190 153776 114246 153785
rect 114190 153711 114246 153720
rect 114098 86864 114154 86873
rect 114098 86799 114154 86808
rect 114204 85377 114232 153711
rect 114282 151056 114338 151065
rect 114282 150991 114338 151000
rect 114190 85368 114246 85377
rect 114190 85303 114246 85312
rect 114296 82385 114324 150991
rect 114388 103193 114416 214639
rect 115846 214568 115902 214577
rect 115846 214503 115902 214512
rect 115754 208992 115810 209001
rect 115754 208927 115810 208936
rect 114466 203552 114522 203561
rect 114466 203487 114522 203496
rect 114374 103184 114430 103193
rect 114374 103119 114430 103128
rect 114376 89684 114428 89690
rect 114376 89626 114428 89632
rect 114282 82376 114338 82385
rect 114282 82311 114338 82320
rect 113822 80880 113878 80889
rect 113822 80815 113878 80824
rect 114388 80186 114416 89626
rect 114480 83745 114508 203487
rect 115662 149696 115718 149705
rect 115662 149631 115718 149640
rect 115478 141400 115534 141409
rect 115478 141335 115534 141344
rect 115386 136096 115442 136105
rect 115386 136031 115442 136040
rect 115400 101833 115428 136031
rect 115386 101824 115442 101833
rect 115386 101759 115442 101768
rect 115492 98841 115520 141335
rect 115570 135960 115626 135969
rect 115570 135895 115626 135904
rect 115478 98832 115534 98841
rect 115478 98767 115534 98776
rect 115584 92449 115612 135895
rect 115676 95237 115704 149631
rect 115768 96733 115796 208927
rect 115754 96724 115810 96733
rect 115754 96659 115810 96668
rect 115662 95228 115718 95237
rect 115662 95163 115718 95172
rect 115860 93741 115888 214503
rect 116766 195256 116822 195265
rect 116766 195191 116822 195200
rect 116584 180736 116636 180742
rect 116584 180678 116636 180684
rect 116492 129872 116544 129878
rect 116490 129840 116492 129849
rect 116544 129840 116546 129849
rect 116490 129775 116546 129784
rect 116492 100360 116544 100366
rect 116490 100328 116492 100337
rect 116544 100328 116546 100337
rect 116490 100263 116546 100272
rect 115846 93732 115902 93741
rect 115846 93667 115902 93676
rect 115570 92440 115626 92449
rect 115570 92375 115626 92384
rect 114466 83736 114522 83745
rect 114466 83671 114522 83680
rect 114388 80158 114600 80186
rect 114374 76664 114430 76673
rect 114374 76599 114430 76608
rect 112536 74384 112588 74390
rect 112536 74326 112588 74332
rect 112444 74248 112496 74254
rect 112444 74190 112496 74196
rect 113916 72820 113968 72826
rect 113916 72762 113968 72768
rect 109684 72684 109736 72690
rect 109684 72626 109736 72632
rect 107016 72548 107068 72554
rect 107016 72490 107068 72496
rect 105726 71224 105782 71233
rect 105726 71159 105782 71168
rect 104162 70136 104218 70145
rect 104162 70071 104218 70080
rect 90362 69728 90418 69737
rect 90362 69663 90418 69672
rect 86868 65748 86920 65754
rect 86868 65690 86920 65696
rect 85672 13116 85724 13122
rect 85672 13058 85724 13064
rect 85684 480 85712 13058
rect 86880 480 86908 65690
rect 87970 61432 88026 61441
rect 87970 61367 88026 61376
rect 87984 480 88012 61367
rect 89166 6216 89222 6225
rect 89166 6151 89222 6160
rect 89180 480 89208 6151
rect 90376 480 90404 69663
rect 105544 68604 105596 68610
rect 105544 68546 105596 68552
rect 93952 68536 94004 68542
rect 93952 68478 94004 68484
rect 91558 55856 91614 55865
rect 91558 55791 91614 55800
rect 91572 480 91600 55791
rect 92756 47660 92808 47666
rect 92756 47602 92808 47608
rect 92768 480 92796 47602
rect 93964 480 93992 68478
rect 103336 67108 103388 67114
rect 103336 67050 103388 67056
rect 97448 67040 97500 67046
rect 97448 66982 97500 66988
rect 95148 44940 95200 44946
rect 95148 44882 95200 44888
rect 95160 480 95188 44882
rect 96252 8968 96304 8974
rect 96252 8910 96304 8916
rect 96264 480 96292 8910
rect 97460 480 97488 66982
rect 101036 65816 101088 65822
rect 101036 65758 101088 65764
rect 99840 49020 99892 49026
rect 99840 48962 99892 48968
rect 98644 3800 98696 3806
rect 98644 3742 98696 3748
rect 98656 480 98684 3742
rect 99852 480 99880 48962
rect 101048 480 101076 65758
rect 102232 62960 102284 62966
rect 102232 62902 102284 62908
rect 102244 480 102272 62902
rect 103348 480 103376 67050
rect 105556 3262 105584 68546
rect 104532 3256 104584 3262
rect 104532 3198 104584 3204
rect 105544 3256 105596 3262
rect 105544 3198 105596 3204
rect 104544 480 104572 3198
rect 105740 480 105768 71159
rect 106924 57384 106976 57390
rect 106924 57326 106976 57332
rect 106936 480 106964 57326
rect 107028 25566 107056 72490
rect 109316 61532 109368 61538
rect 109316 61474 109368 61480
rect 107016 25560 107068 25566
rect 107016 25502 107068 25508
rect 108120 3868 108172 3874
rect 108120 3810 108172 3816
rect 108132 480 108160 3810
rect 109328 480 109356 61474
rect 109696 17270 109724 72626
rect 111064 71256 111116 71262
rect 111064 71198 111116 71204
rect 109684 17264 109736 17270
rect 109684 17206 109736 17212
rect 111076 3806 111104 71198
rect 113824 68672 113876 68678
rect 113824 68614 113876 68620
rect 112444 65884 112496 65890
rect 112444 65826 112496 65832
rect 111064 3800 111116 3806
rect 111064 3742 111116 3748
rect 112456 3398 112484 65826
rect 112812 64388 112864 64394
rect 112812 64330 112864 64336
rect 110512 3392 110564 3398
rect 110512 3334 110564 3340
rect 112444 3392 112496 3398
rect 112444 3334 112496 3340
rect 110524 480 110552 3334
rect 111616 3256 111668 3262
rect 111616 3198 111668 3204
rect 111628 480 111656 3198
rect 112824 480 112852 64330
rect 113836 3262 113864 68614
rect 113928 15910 113956 72762
rect 114388 59673 114416 76599
rect 114572 75682 114600 80158
rect 116490 78160 116546 78169
rect 116490 78095 116546 78104
rect 114560 75676 114612 75682
rect 114560 75618 114612 75624
rect 116504 75585 116532 78095
rect 116490 75576 116546 75585
rect 116490 75511 116546 75520
rect 114466 75168 114522 75177
rect 114466 75103 114522 75112
rect 114374 59664 114430 59673
rect 114374 59599 114430 59608
rect 114480 58585 114508 75103
rect 116400 70780 116452 70786
rect 116400 70722 116452 70728
rect 115204 67176 115256 67182
rect 115204 67118 115256 67124
rect 114466 58576 114522 58585
rect 114466 58511 114522 58520
rect 114008 58404 114060 58410
rect 114008 58346 114060 58352
rect 113916 15904 113968 15910
rect 113916 15846 113968 15852
rect 113824 3256 113876 3262
rect 113824 3198 113876 3204
rect 114020 480 114048 58346
rect 115216 480 115244 67118
rect 116412 480 116440 70722
rect 116596 69494 116624 180678
rect 116674 139360 116730 139369
rect 116674 139295 116730 139304
rect 116688 129878 116716 139295
rect 116676 129872 116728 129878
rect 116676 129814 116728 129820
rect 116780 100366 116808 195191
rect 117240 180713 117268 214540
rect 146312 214526 146510 214554
rect 146312 207097 146340 214526
rect 149072 213217 149100 215863
rect 396460 214849 396488 285631
rect 177854 214840 177910 214849
rect 177854 214775 177910 214784
rect 390558 214840 390614 214849
rect 390558 214775 390614 214784
rect 396446 214840 396502 214849
rect 396446 214775 396502 214784
rect 149058 213208 149114 213217
rect 149058 213143 149114 213152
rect 159362 213208 159418 213217
rect 159362 213143 159418 213152
rect 162122 213208 162178 213217
rect 162122 213143 162178 213152
rect 159376 209137 159404 213143
rect 159362 209128 159418 209137
rect 159362 209063 159418 209072
rect 143446 207088 143502 207097
rect 143446 207023 143502 207032
rect 146298 207088 146354 207097
rect 146298 207023 146354 207032
rect 134522 193896 134578 193905
rect 134522 193831 134578 193840
rect 134536 184006 134564 193831
rect 134524 184000 134576 184006
rect 134524 183942 134576 183948
rect 137284 184000 137336 184006
rect 143460 183954 143488 207023
rect 149520 191140 149572 191146
rect 149520 191082 149572 191088
rect 147588 189780 147640 189786
rect 147588 189722 147640 189728
rect 146208 188352 146260 188358
rect 146208 188294 146260 188300
rect 144736 185632 144788 185638
rect 144736 185574 144788 185580
rect 137336 183948 137586 183954
rect 137284 183942 137586 183948
rect 137296 183926 137586 183942
rect 143198 183926 143488 183954
rect 144748 183940 144776 185574
rect 146220 183940 146248 188294
rect 147600 183940 147628 189722
rect 149532 183940 149560 191082
rect 157246 186960 157302 186969
rect 157246 186895 157302 186904
rect 152738 184240 152794 184249
rect 152738 184175 152794 184184
rect 152752 183940 152780 184175
rect 155958 183560 156014 183569
rect 155958 183495 156014 183504
rect 157260 183433 157288 186895
rect 154302 183424 154358 183433
rect 154302 183359 154358 183368
rect 157246 183424 157302 183433
rect 157246 183359 157302 183368
rect 151202 182566 151584 182594
rect 151556 182510 151584 182566
rect 151544 182504 151596 182510
rect 151544 182446 151596 182452
rect 154488 182504 154540 182510
rect 154488 182446 154540 182452
rect 138572 182436 138624 182442
rect 138572 182378 138624 182384
rect 133234 182064 133290 182073
rect 133234 181999 133236 182008
rect 133288 181999 133290 182008
rect 136638 182064 136694 182073
rect 136638 181999 136640 182008
rect 133236 181970 133288 181976
rect 136692 181999 136694 182008
rect 136640 181970 136692 181976
rect 136548 181552 136600 181558
rect 136548 181494 136600 181500
rect 118608 181212 118660 181218
rect 118608 181154 118660 181160
rect 117226 180704 117282 180713
rect 117226 180639 117282 180648
rect 118620 142154 118648 181154
rect 128268 181008 128320 181014
rect 128268 180950 128320 180956
rect 120724 178696 120776 178702
rect 120724 178638 120776 178644
rect 118160 142126 118648 142154
rect 118160 134994 118188 142126
rect 120736 137018 120764 178638
rect 121368 177336 121420 177342
rect 121368 177278 121420 177284
rect 121380 142154 121408 177278
rect 124864 175908 124916 175914
rect 124864 175850 124916 175856
rect 121288 142126 121408 142154
rect 119344 137012 119396 137018
rect 119344 136954 119396 136960
rect 120724 137012 120776 137018
rect 120724 136954 120776 136960
rect 117806 134966 118188 134994
rect 119356 134980 119384 136954
rect 121288 134994 121316 142126
rect 124876 137970 124904 175850
rect 128280 142154 128308 180950
rect 133234 180704 133290 180713
rect 133234 180639 133290 180648
rect 129648 179512 129700 179518
rect 129648 179454 129700 179460
rect 129660 142154 129688 179454
rect 133248 179450 133276 180639
rect 136364 179512 136416 179518
rect 136362 179480 136364 179489
rect 136416 179480 136418 179489
rect 133236 179444 133288 179450
rect 136362 179415 136418 179424
rect 133236 179386 133288 179392
rect 136560 178702 136588 181494
rect 138584 181393 138612 182378
rect 146024 181620 146076 181626
rect 146024 181562 146076 181568
rect 138570 181384 138626 181393
rect 138570 181319 138626 181328
rect 137834 181248 137890 181257
rect 138754 181248 138810 181257
rect 138032 181218 138138 181234
rect 137834 181183 137890 181192
rect 138020 181212 138138 181218
rect 137848 181150 137876 181183
rect 138072 181206 138138 181212
rect 138676 181206 138754 181234
rect 138020 181154 138072 181160
rect 137836 181144 137888 181150
rect 137836 181086 137888 181092
rect 137928 181144 137980 181150
rect 137928 181086 137980 181092
rect 138018 181112 138074 181121
rect 136548 178696 136600 178702
rect 136548 178638 136600 178644
rect 137940 177342 137968 181086
rect 138676 181084 138704 181206
rect 138754 181183 138810 181192
rect 138018 181047 138020 181056
rect 138072 181047 138074 181056
rect 138020 181018 138072 181024
rect 146036 180878 146064 181562
rect 154500 181393 154528 182446
rect 154672 182436 154724 182442
rect 154672 182378 154724 182384
rect 154486 181384 154542 181393
rect 154486 181319 154542 181328
rect 146024 180872 146076 180878
rect 146024 180814 146076 180820
rect 146024 180600 146076 180606
rect 146024 180542 146076 180548
rect 140962 179752 141018 179761
rect 140962 179687 141018 179696
rect 140976 179450 141004 179687
rect 146036 179625 146064 180542
rect 149886 180024 149942 180033
rect 149886 179959 149942 179968
rect 146022 179616 146078 179625
rect 146022 179551 146078 179560
rect 146298 179480 146354 179489
rect 140964 179444 141016 179450
rect 146298 179415 146354 179424
rect 140964 179386 141016 179392
rect 137928 177336 137980 177342
rect 137928 177278 137980 177284
rect 146312 177070 146340 179415
rect 149900 177970 149928 179959
rect 151726 179888 151782 179897
rect 151726 179823 151782 179832
rect 150990 179752 151046 179761
rect 150990 179687 151046 179696
rect 151004 177970 151032 179687
rect 149638 177942 149928 177970
rect 150742 177942 151032 177970
rect 151740 177820 151768 179823
rect 154684 177818 154712 182378
rect 162136 181801 162164 213143
rect 176672 211138 176700 214540
rect 176842 211848 176898 211857
rect 176842 211783 176898 211792
rect 174544 211132 174596 211138
rect 174544 211074 174596 211080
rect 176660 211132 176712 211138
rect 176660 211074 176712 211080
rect 167642 209128 167698 209137
rect 167642 209063 167698 209072
rect 167656 198801 167684 209063
rect 167642 198792 167698 198801
rect 167642 198727 167698 198736
rect 173162 198792 173218 198801
rect 173162 198727 173218 198736
rect 173176 186425 173204 198727
rect 173162 186416 173218 186425
rect 173162 186351 173218 186360
rect 174556 185638 174584 211074
rect 175278 210352 175334 210361
rect 175278 210287 175334 210296
rect 174544 185632 174596 185638
rect 174544 185574 174596 185580
rect 155774 181792 155830 181801
rect 155774 181727 155830 181736
rect 162122 181792 162178 181801
rect 162122 181727 162178 181736
rect 155406 181384 155462 181393
rect 155788 181370 155816 181727
rect 155462 181342 155816 181370
rect 163042 181384 163098 181393
rect 155406 181319 155462 181328
rect 163042 181319 163098 181328
rect 155500 180532 155552 180538
rect 155500 180474 155552 180480
rect 161480 180532 161532 180538
rect 161480 180474 161532 180480
rect 155408 180396 155460 180402
rect 155408 180338 155460 180344
rect 155420 180033 155448 180338
rect 155406 180024 155462 180033
rect 155406 179959 155462 179968
rect 155512 179897 155540 180474
rect 155776 180464 155828 180470
rect 155776 180406 155828 180412
rect 155498 179888 155554 179897
rect 155498 179823 155554 179832
rect 155788 179761 155816 180406
rect 155774 179752 155830 179761
rect 155774 179687 155830 179696
rect 154672 177812 154724 177818
rect 154672 177754 154724 177760
rect 141516 177064 141568 177070
rect 141358 177012 141516 177018
rect 141358 177006 141568 177012
rect 146300 177064 146352 177070
rect 146300 177006 146352 177012
rect 141358 176990 141556 177006
rect 161492 176526 161520 180474
rect 162766 179480 162822 179489
rect 162766 179415 162822 179424
rect 162780 177886 162808 179415
rect 162768 177880 162820 177886
rect 162768 177822 162820 177828
rect 161480 176520 161532 176526
rect 161480 176462 161532 176468
rect 163056 176460 163084 181319
rect 163504 180464 163556 180470
rect 163504 180406 163556 180412
rect 142618 176080 142674 176089
rect 138584 175914 138612 175916
rect 138572 175908 138624 175914
rect 138572 175850 138624 175856
rect 141896 172553 141924 176052
rect 142674 176038 142922 176066
rect 142618 176015 142674 176024
rect 161480 175908 161532 175914
rect 161480 175850 161532 175856
rect 161492 175386 161520 175850
rect 161400 175358 161520 175386
rect 161400 175030 161428 175358
rect 161388 175024 161440 175030
rect 161388 174966 161440 174972
rect 161388 174752 161440 174758
rect 161388 174694 161440 174700
rect 161400 174298 161428 174694
rect 161400 174270 161520 174298
rect 141882 172544 141938 172553
rect 141882 172479 141938 172488
rect 161492 167618 161520 174270
rect 161480 167612 161532 167618
rect 161480 167554 161532 167560
rect 161480 167340 161532 167346
rect 161480 167282 161532 167288
rect 139490 165200 139546 165209
rect 139490 165135 139546 165144
rect 136086 162072 136142 162081
rect 136362 162072 136418 162081
rect 136142 162030 136362 162058
rect 136086 162007 136142 162016
rect 136362 162007 136418 162016
rect 137848 161498 137954 161514
rect 136456 161492 136508 161498
rect 136456 161434 136508 161440
rect 137836 161492 137954 161498
rect 137888 161486 137954 161492
rect 137836 161434 137888 161440
rect 136468 161226 136496 161434
rect 135444 161220 135496 161226
rect 135444 161162 135496 161168
rect 136456 161220 136508 161226
rect 136456 161162 136508 161168
rect 133788 158772 133840 158778
rect 133788 158714 133840 158720
rect 132408 158092 132460 158098
rect 132408 158034 132460 158040
rect 131028 157412 131080 157418
rect 131028 157354 131080 157360
rect 131040 142154 131068 157354
rect 132420 142154 132448 158034
rect 127544 142126 128308 142154
rect 129200 142126 129688 142154
rect 130672 142126 131068 142154
rect 132328 142126 132448 142154
rect 124036 137964 124088 137970
rect 124036 137906 124088 137912
rect 124864 137964 124916 137970
rect 124864 137906 124916 137912
rect 122470 137456 122526 137465
rect 122470 137391 122526 137400
rect 120934 134966 121316 134994
rect 122484 134980 122512 137391
rect 124048 134980 124076 137906
rect 125598 137592 125654 137601
rect 125598 137527 125654 137536
rect 125612 134980 125640 137527
rect 127544 134994 127572 142126
rect 129200 134994 129228 142126
rect 130672 134994 130700 142126
rect 132328 134994 132356 142126
rect 133800 134994 133828 158714
rect 134536 157418 134564 159732
rect 134524 157412 134576 157418
rect 134524 157354 134576 157360
rect 135456 151814 135484 161162
rect 139504 161129 139532 165135
rect 147496 162648 147548 162654
rect 147496 162590 147548 162596
rect 147508 162588 147536 162590
rect 161492 161770 161520 167282
rect 161480 161764 161532 161770
rect 161480 161706 161532 161712
rect 163228 161628 163280 161634
rect 163228 161570 163280 161576
rect 163240 161537 163268 161570
rect 160466 161528 160522 161537
rect 163226 161528 163282 161537
rect 160466 161463 160468 161472
rect 160520 161463 160522 161472
rect 161480 161492 161532 161498
rect 160468 161434 160520 161440
rect 163226 161463 163282 161472
rect 161480 161434 161532 161440
rect 139490 161120 139546 161129
rect 139490 161055 139546 161064
rect 135640 158098 135668 159732
rect 136652 158778 136680 159732
rect 136640 158772 136692 158778
rect 136640 158714 136692 158720
rect 135628 158092 135680 158098
rect 135628 158034 135680 158040
rect 138676 157418 138704 159732
rect 139688 157434 139716 159732
rect 140792 157434 140820 159732
rect 136548 157412 136600 157418
rect 136548 157354 136600 157360
rect 138664 157412 138716 157418
rect 138664 157354 138716 157360
rect 139320 157406 139716 157434
rect 140700 157406 140820 157434
rect 135456 151786 136496 151814
rect 136468 137902 136496 151786
rect 134984 137896 135036 137902
rect 134984 137838 135036 137844
rect 136456 137896 136508 137902
rect 136456 137838 136508 137844
rect 127190 134966 127572 134994
rect 128754 134966 129228 134994
rect 130318 134966 130700 134994
rect 131882 134966 132356 134994
rect 133446 134966 133828 134994
rect 134996 134980 135024 137838
rect 136560 134980 136588 157354
rect 139320 142154 139348 157406
rect 140700 142154 140728 157406
rect 141620 142154 141648 159732
rect 138584 142126 139348 142154
rect 140056 142126 140728 142154
rect 141436 142126 141648 142154
rect 138584 134994 138612 142126
rect 140056 134994 140084 142126
rect 141436 134994 141464 142126
rect 138138 134966 138612 134994
rect 139702 134966 140084 134994
rect 141266 134966 141464 134994
rect 142816 134980 142844 159732
rect 144196 134994 144224 159732
rect 145406 159718 145512 159746
rect 145484 151814 145512 159718
rect 145484 151786 145604 151814
rect 145576 134994 145604 151786
rect 146220 137970 146248 159732
rect 147338 159718 147536 159746
rect 148350 159718 148548 159746
rect 147508 151814 147536 159718
rect 148520 155786 148548 159718
rect 148508 155780 148560 155786
rect 148508 155722 148560 155728
rect 147508 151786 147628 151814
rect 146208 137964 146260 137970
rect 146208 137906 146260 137912
rect 147496 137964 147548 137970
rect 147496 137906 147548 137912
rect 144196 134966 144394 134994
rect 145576 134966 145958 134994
rect 147508 134980 147536 137906
rect 147600 136814 147628 151786
rect 148888 137834 148916 159732
rect 148968 155780 149020 155786
rect 148968 155722 149020 155728
rect 148876 137828 148928 137834
rect 148876 137770 148928 137776
rect 148980 137018 149008 155722
rect 150360 137902 150388 159732
rect 151372 157418 151400 159732
rect 151360 157412 151412 157418
rect 151360 157354 151412 157360
rect 152464 157412 152516 157418
rect 152464 157354 152516 157360
rect 152476 137970 152504 157354
rect 152464 137964 152516 137970
rect 152464 137906 152516 137912
rect 155316 137964 155368 137970
rect 155316 137906 155368 137912
rect 150348 137896 150400 137902
rect 150348 137838 150400 137844
rect 153752 137896 153804 137902
rect 153752 137838 153804 137844
rect 152188 137828 152240 137834
rect 152188 137770 152240 137776
rect 148968 137012 149020 137018
rect 148968 136954 149020 136960
rect 150624 137012 150676 137018
rect 150624 136954 150676 136960
rect 147588 136808 147640 136814
rect 147588 136750 147640 136756
rect 149060 136808 149112 136814
rect 149060 136750 149112 136756
rect 149072 134980 149100 136750
rect 150636 134980 150664 136954
rect 152200 134980 152228 137770
rect 153764 134980 153792 137838
rect 155328 134980 155356 137906
rect 156880 137692 156932 137698
rect 156880 137634 156932 137640
rect 156892 134980 156920 137634
rect 161400 137358 161428 159732
rect 161388 137352 161440 137358
rect 161388 137294 161440 137300
rect 158444 137148 158496 137154
rect 158444 137090 158496 137096
rect 158456 134980 158484 137090
rect 161492 136746 161520 161434
rect 162334 159718 162532 159746
rect 161570 152416 161626 152425
rect 161570 152351 161626 152360
rect 160008 136740 160060 136746
rect 160008 136682 160060 136688
rect 161480 136740 161532 136746
rect 161480 136682 161532 136688
rect 160020 134980 160048 136682
rect 161584 134980 161612 152351
rect 162504 151814 162532 159718
rect 163332 159390 163360 159732
rect 163320 159384 163372 159390
rect 163320 159326 163372 159332
rect 162504 151786 162808 151814
rect 162780 137290 162808 151786
rect 162768 137284 162820 137290
rect 162768 137226 162820 137232
rect 163516 137154 163544 180406
rect 163596 180396 163648 180402
rect 163596 180338 163648 180344
rect 163608 137698 163636 180338
rect 164884 177880 164936 177886
rect 164884 177822 164936 177828
rect 164240 161628 164292 161634
rect 164240 161570 164292 161576
rect 163686 160712 163742 160721
rect 163686 160647 163742 160656
rect 163596 137692 163648 137698
rect 163596 137634 163648 137640
rect 163504 137148 163556 137154
rect 163504 137090 163556 137096
rect 163700 134994 163728 160647
rect 163162 134966 163728 134994
rect 164252 134994 164280 161570
rect 164896 146266 164924 177822
rect 168378 162208 168434 162217
rect 168378 162143 168434 162152
rect 168392 151814 168420 162143
rect 173900 159384 173952 159390
rect 173900 159326 173952 159332
rect 168392 151786 169064 151814
rect 164884 146260 164936 146266
rect 164884 146202 164936 146208
rect 165896 146260 165948 146266
rect 165896 146202 165948 146208
rect 165908 134994 165936 146202
rect 167826 137456 167882 137465
rect 167826 137391 167882 137400
rect 164252 134966 164726 134994
rect 165908 134966 166290 134994
rect 167840 134980 167868 137391
rect 169036 134994 169064 151786
rect 170956 137352 171008 137358
rect 170956 137294 171008 137300
rect 169036 134966 169418 134994
rect 170968 134980 170996 137294
rect 172520 137284 172572 137290
rect 172520 137226 172572 137232
rect 172532 134980 172560 137226
rect 173912 134994 173940 159326
rect 175292 151814 175320 210287
rect 175922 186416 175978 186425
rect 175922 186351 175978 186360
rect 175292 151786 175412 151814
rect 173912 134966 174110 134994
rect 175384 126993 175412 151786
rect 175370 126984 175426 126993
rect 175370 126919 175426 126928
rect 175936 118833 175964 186351
rect 176750 162072 176806 162081
rect 176750 162007 176806 162016
rect 176658 134464 176714 134473
rect 176658 134399 176714 134408
rect 175922 118824 175978 118833
rect 175922 118759 175978 118768
rect 176672 107545 176700 134399
rect 176764 128353 176792 162007
rect 176750 128344 176806 128353
rect 176750 128279 176806 128288
rect 176856 125497 176884 211783
rect 177304 210452 177356 210458
rect 177304 210394 177356 210400
rect 176934 141536 176990 141545
rect 176934 141471 176990 141480
rect 176842 125488 176898 125497
rect 176842 125423 176898 125432
rect 176948 111761 176976 141471
rect 177026 132560 177082 132569
rect 177026 132495 177082 132504
rect 176934 111752 176990 111761
rect 176934 111687 176990 111696
rect 176658 107536 176714 107545
rect 176658 107471 176714 107480
rect 116768 100360 116820 100366
rect 116768 100302 116820 100308
rect 116676 84244 116728 84250
rect 116676 84186 116728 84192
rect 116688 74322 116716 84186
rect 175280 76560 175332 76566
rect 175280 76502 175332 76508
rect 119988 75676 120040 75682
rect 119988 75618 120040 75624
rect 170496 75676 170548 75682
rect 170496 75618 170548 75624
rect 170588 75676 170640 75682
rect 170588 75618 170640 75624
rect 170680 75676 170732 75682
rect 170680 75618 170732 75624
rect 120000 74474 120028 75618
rect 170404 75540 170456 75546
rect 170404 75482 170456 75488
rect 121472 75126 121578 75154
rect 120000 74446 120120 74474
rect 116676 74316 116728 74322
rect 116676 74258 116728 74264
rect 117870 73128 117926 73137
rect 117870 73063 117926 73072
rect 119620 73092 119672 73098
rect 117884 72593 117912 73063
rect 119620 73034 119672 73040
rect 118148 72752 118200 72758
rect 118148 72694 118200 72700
rect 117870 72584 117926 72593
rect 117870 72519 117926 72528
rect 116858 72040 116914 72049
rect 116858 71975 116914 71984
rect 116768 71868 116820 71874
rect 116768 71810 116820 71816
rect 116674 69592 116730 69601
rect 116674 69527 116730 69536
rect 116584 69488 116636 69494
rect 116584 69430 116636 69436
rect 116688 3534 116716 69527
rect 116780 7614 116808 71810
rect 116872 18630 116900 71975
rect 118056 71800 118108 71806
rect 118056 71742 118108 71748
rect 117964 71596 118016 71602
rect 117964 71538 118016 71544
rect 117976 71126 118004 71538
rect 117964 71120 118016 71126
rect 117964 71062 118016 71068
rect 117962 70408 118018 70417
rect 117962 70343 118018 70352
rect 117596 68740 117648 68746
rect 117596 68682 117648 68688
rect 117228 60852 117280 60858
rect 117228 60794 117280 60800
rect 117240 60042 117268 60794
rect 117228 60036 117280 60042
rect 117228 59978 117280 59984
rect 116860 18624 116912 18630
rect 116860 18566 116912 18572
rect 116768 7608 116820 7614
rect 116768 7550 116820 7556
rect 116676 3528 116728 3534
rect 116676 3470 116728 3476
rect 117608 480 117636 68682
rect 117976 3466 118004 70343
rect 118068 10334 118096 71742
rect 118160 14482 118188 72694
rect 119344 72072 119396 72078
rect 119344 72014 119396 72020
rect 118792 70032 118844 70038
rect 118792 69974 118844 69980
rect 118148 14476 118200 14482
rect 118148 14418 118200 14424
rect 118056 10328 118108 10334
rect 118056 10270 118108 10276
rect 117964 3460 118016 3466
rect 117964 3402 118016 3408
rect 118804 480 118832 69974
rect 119356 3874 119384 72014
rect 119436 71732 119488 71738
rect 119436 71674 119488 71680
rect 119344 3868 119396 3874
rect 119344 3810 119396 3816
rect 119448 3602 119476 71674
rect 119528 69080 119580 69086
rect 119528 69022 119580 69028
rect 119540 3670 119568 69022
rect 119632 58410 119660 73034
rect 120092 71777 120120 74446
rect 121184 73024 121236 73030
rect 120262 72992 120318 73001
rect 121184 72966 121236 72972
rect 120262 72927 120318 72936
rect 120276 72729 120304 72927
rect 120262 72720 120318 72729
rect 120262 72655 120318 72664
rect 121000 72344 121052 72350
rect 121000 72286 121052 72292
rect 120908 72276 120960 72282
rect 120908 72218 120960 72224
rect 120724 71936 120776 71942
rect 120724 71878 120776 71884
rect 120078 71768 120134 71777
rect 120078 71703 120134 71712
rect 119620 58404 119672 58410
rect 119620 58346 119672 58352
rect 120736 4894 120764 71878
rect 120816 71664 120868 71670
rect 120816 71606 120868 71612
rect 120724 4888 120776 4894
rect 120724 4830 120776 4836
rect 120828 3738 120856 71606
rect 120920 13122 120948 72218
rect 121012 40730 121040 72286
rect 121092 71324 121144 71330
rect 121092 71266 121144 71272
rect 121000 40724 121052 40730
rect 121000 40666 121052 40672
rect 120908 13116 120960 13122
rect 120908 13058 120960 13064
rect 120816 3732 120868 3738
rect 120816 3674 120868 3680
rect 119528 3664 119580 3670
rect 119528 3606 119580 3612
rect 119436 3596 119488 3602
rect 119436 3538 119488 3544
rect 119896 3460 119948 3466
rect 119896 3402 119948 3408
rect 119908 480 119936 3402
rect 121104 480 121132 71266
rect 121196 49026 121224 72966
rect 121276 72820 121328 72826
rect 121276 72762 121328 72768
rect 121288 57390 121316 72762
rect 121472 70553 121500 75126
rect 121656 72729 121684 75140
rect 121642 72720 121698 72729
rect 121642 72655 121698 72664
rect 121458 70544 121514 70553
rect 121748 70530 121776 75140
rect 121458 70479 121514 70488
rect 121656 70502 121776 70530
rect 121552 65952 121604 65958
rect 121552 65894 121604 65900
rect 121564 65754 121592 65894
rect 121552 65748 121604 65754
rect 121552 65690 121604 65696
rect 121656 65550 121684 70502
rect 121736 70440 121788 70446
rect 121736 70382 121788 70388
rect 121748 68338 121776 70382
rect 121736 68332 121788 68338
rect 121736 68274 121788 68280
rect 121840 65686 121868 75140
rect 121932 73001 121960 75140
rect 121918 72992 121974 73001
rect 121918 72927 121974 72936
rect 122024 67634 122052 75140
rect 122116 70446 122144 75140
rect 122104 70440 122156 70446
rect 122104 70382 122156 70388
rect 122024 67606 122144 67634
rect 121920 66020 121972 66026
rect 121920 65962 121972 65968
rect 121828 65680 121880 65686
rect 121828 65622 121880 65628
rect 121644 65544 121696 65550
rect 121644 65486 121696 65492
rect 121736 65544 121788 65550
rect 121736 65486 121788 65492
rect 121276 57384 121328 57390
rect 121276 57326 121328 57332
rect 121748 51746 121776 65486
rect 121932 65226 121960 65962
rect 121840 65198 121960 65226
rect 121840 57254 121868 65198
rect 122116 57974 122144 67606
rect 122208 66026 122236 75140
rect 122196 66020 122248 66026
rect 122196 65962 122248 65968
rect 122300 60858 122328 75140
rect 122392 72049 122420 75140
rect 122378 72040 122434 72049
rect 122378 71975 122434 71984
rect 122380 65680 122432 65686
rect 122380 65622 122432 65628
rect 122288 60852 122340 60858
rect 122288 60794 122340 60800
rect 122392 60734 122420 65622
rect 122484 64190 122512 75140
rect 122576 65550 122604 75140
rect 122564 65544 122616 65550
rect 122564 65486 122616 65492
rect 122472 64184 122524 64190
rect 122472 64126 122524 64132
rect 122300 60706 122420 60734
rect 122116 57946 122236 57974
rect 121828 57248 121880 57254
rect 121828 57190 121880 57196
rect 121736 51740 121788 51746
rect 121736 51682 121788 51688
rect 121184 49020 121236 49026
rect 121184 48962 121236 48968
rect 122208 6186 122236 57946
rect 122300 46238 122328 60706
rect 122668 50386 122696 75140
rect 122760 71738 122788 75140
rect 122852 72457 122880 75140
rect 122944 73370 122972 75140
rect 122932 73364 122984 73370
rect 122932 73306 122984 73312
rect 123036 73250 123064 75140
rect 122944 73222 123064 73250
rect 122838 72448 122894 72457
rect 122838 72383 122894 72392
rect 122840 72004 122892 72010
rect 122840 71946 122892 71952
rect 122748 71732 122800 71738
rect 122748 71674 122800 71680
rect 122656 50380 122708 50386
rect 122656 50322 122708 50328
rect 122288 46232 122340 46238
rect 122288 46174 122340 46180
rect 122852 16574 122880 71946
rect 122944 71806 122972 73222
rect 123128 73114 123156 75140
rect 123036 73086 123156 73114
rect 123036 72554 123064 73086
rect 123116 72956 123168 72962
rect 123116 72898 123168 72904
rect 123024 72548 123076 72554
rect 123024 72490 123076 72496
rect 122932 71800 122984 71806
rect 122932 71742 122984 71748
rect 123128 65618 123156 72898
rect 123220 72729 123248 75140
rect 123206 72720 123262 72729
rect 123206 72655 123262 72664
rect 123208 72616 123260 72622
rect 123208 72558 123260 72564
rect 123220 71874 123248 72558
rect 123312 72486 123340 75140
rect 123404 72690 123432 75140
rect 123392 72684 123444 72690
rect 123392 72626 123444 72632
rect 123390 72584 123446 72593
rect 123390 72519 123446 72528
rect 123404 72486 123432 72519
rect 123300 72480 123352 72486
rect 123300 72422 123352 72428
rect 123392 72480 123444 72486
rect 123392 72422 123444 72428
rect 123392 72344 123444 72350
rect 123392 72286 123444 72292
rect 123208 71868 123260 71874
rect 123208 71810 123260 71816
rect 123300 65680 123352 65686
rect 123300 65622 123352 65628
rect 123116 65612 123168 65618
rect 123116 65554 123168 65560
rect 123312 53106 123340 65622
rect 123404 54534 123432 72286
rect 123496 65414 123524 75140
rect 123588 72962 123616 75140
rect 123680 73545 123708 75140
rect 123666 73536 123722 73545
rect 123666 73471 123722 73480
rect 123668 73364 123720 73370
rect 123668 73306 123720 73312
rect 123576 72956 123628 72962
rect 123576 72898 123628 72904
rect 123574 72856 123630 72865
rect 123574 72791 123630 72800
rect 123588 72622 123616 72791
rect 123576 72616 123628 72622
rect 123576 72558 123628 72564
rect 123576 72140 123628 72146
rect 123576 72082 123628 72088
rect 123484 65408 123536 65414
rect 123484 65350 123536 65356
rect 123588 55962 123616 72082
rect 123680 71097 123708 73306
rect 123772 72758 123800 75140
rect 123760 72752 123812 72758
rect 123760 72694 123812 72700
rect 123758 72584 123814 72593
rect 123758 72519 123814 72528
rect 123666 71088 123722 71097
rect 123666 71023 123722 71032
rect 123772 70922 123800 72519
rect 123760 70916 123812 70922
rect 123760 70858 123812 70864
rect 123864 68406 123892 75140
rect 123852 68400 123904 68406
rect 123852 68342 123904 68348
rect 123956 65686 123984 75140
rect 123944 65680 123996 65686
rect 123944 65622 123996 65628
rect 124048 65532 124076 75140
rect 124140 72350 124168 75140
rect 124232 72729 124260 75140
rect 124324 73234 124352 75140
rect 124312 73228 124364 73234
rect 124312 73170 124364 73176
rect 124310 73128 124366 73137
rect 124310 73063 124366 73072
rect 124218 72720 124274 72729
rect 124218 72655 124274 72664
rect 124324 72554 124352 73063
rect 124416 72593 124444 75140
rect 124508 72729 124536 75140
rect 124600 72865 124628 75140
rect 124586 72856 124642 72865
rect 124586 72791 124642 72800
rect 124588 72752 124640 72758
rect 124494 72720 124550 72729
rect 124588 72694 124640 72700
rect 124494 72655 124550 72664
rect 124402 72584 124458 72593
rect 124312 72548 124364 72554
rect 124402 72519 124458 72528
rect 124312 72490 124364 72496
rect 124600 72434 124628 72694
rect 124232 72406 124628 72434
rect 124128 72344 124180 72350
rect 124128 72286 124180 72292
rect 124128 72208 124180 72214
rect 124128 72150 124180 72156
rect 123772 65504 124076 65532
rect 123576 55956 123628 55962
rect 123576 55898 123628 55904
rect 123772 55894 123800 65504
rect 123852 65408 123904 65414
rect 123852 65350 123904 65356
rect 123864 58682 123892 65350
rect 124140 64326 124168 72150
rect 124232 69698 124260 72406
rect 124404 72276 124456 72282
rect 124404 72218 124456 72224
rect 124220 69692 124272 69698
rect 124220 69634 124272 69640
rect 124416 66910 124444 72218
rect 124404 66904 124456 66910
rect 124404 66846 124456 66852
rect 124128 64320 124180 64326
rect 124128 64262 124180 64268
rect 124692 61402 124720 75140
rect 124784 71602 124812 75140
rect 124876 72690 124904 75140
rect 124864 72684 124916 72690
rect 124864 72626 124916 72632
rect 124772 71596 124824 71602
rect 124772 71538 124824 71544
rect 124968 62830 124996 75140
rect 124956 62824 125008 62830
rect 124956 62766 125008 62772
rect 124680 61396 124732 61402
rect 124680 61338 124732 61344
rect 125060 60734 125088 75140
rect 125152 65550 125180 75140
rect 125244 72894 125272 75140
rect 125232 72888 125284 72894
rect 125232 72830 125284 72836
rect 125232 72752 125284 72758
rect 125232 72694 125284 72700
rect 125244 69086 125272 72694
rect 125232 69080 125284 69086
rect 125232 69022 125284 69028
rect 125140 65544 125192 65550
rect 125140 65486 125192 65492
rect 125336 64258 125364 75140
rect 125324 64252 125376 64258
rect 125324 64194 125376 64200
rect 125060 60706 125272 60734
rect 123852 58676 123904 58682
rect 123852 58618 123904 58624
rect 123760 55888 123812 55894
rect 123760 55830 123812 55836
rect 123392 54528 123444 54534
rect 123392 54470 123444 54476
rect 123300 53100 123352 53106
rect 123300 53042 123352 53048
rect 122852 16546 123064 16574
rect 122196 6180 122248 6186
rect 122196 6122 122248 6128
rect 122288 6180 122340 6186
rect 122288 6122 122340 6128
rect 122300 480 122328 6122
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 125244 4826 125272 60706
rect 125428 7682 125456 75140
rect 125520 72758 125548 75140
rect 125508 72752 125560 72758
rect 125612 72729 125640 75140
rect 125704 72865 125732 75140
rect 125690 72856 125746 72865
rect 125690 72791 125746 72800
rect 125508 72694 125560 72700
rect 125598 72720 125654 72729
rect 125598 72655 125654 72664
rect 125796 69766 125824 75140
rect 125784 69760 125836 69766
rect 125784 69702 125836 69708
rect 125508 65544 125560 65550
rect 125508 65486 125560 65492
rect 125520 10402 125548 65486
rect 125888 62898 125916 75140
rect 125980 72146 126008 75140
rect 125968 72140 126020 72146
rect 125968 72082 126020 72088
rect 126072 68474 126100 75140
rect 126060 68468 126112 68474
rect 126060 68410 126112 68416
rect 126164 65550 126192 75140
rect 126256 72282 126284 75140
rect 126244 72276 126296 72282
rect 126244 72218 126296 72224
rect 126152 65544 126204 65550
rect 126152 65486 126204 65492
rect 125876 62892 125928 62898
rect 125876 62834 125928 62840
rect 126244 60036 126296 60042
rect 126244 59978 126296 59984
rect 125508 10396 125560 10402
rect 125508 10338 125560 10344
rect 125416 7676 125468 7682
rect 125416 7618 125468 7624
rect 125232 4820 125284 4826
rect 125232 4762 125284 4768
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 124680 2984 124732 2990
rect 124680 2926 124732 2932
rect 124692 480 124720 2926
rect 125888 480 125916 3470
rect 126256 3466 126284 59978
rect 126348 53174 126376 75140
rect 126440 72758 126468 75140
rect 126428 72752 126480 72758
rect 126428 72694 126480 72700
rect 126426 72584 126482 72593
rect 126426 72519 126482 72528
rect 126440 71670 126468 72519
rect 126428 71664 126480 71670
rect 126428 71606 126480 71612
rect 126336 53168 126388 53174
rect 126336 53110 126388 53116
rect 126532 44878 126560 75140
rect 126624 70394 126652 75140
rect 126716 73001 126744 75140
rect 126702 72992 126758 73001
rect 126702 72927 126758 72936
rect 126808 72842 126836 75140
rect 126716 72814 126836 72842
rect 126716 72214 126744 72814
rect 126796 72752 126848 72758
rect 126796 72694 126848 72700
rect 126704 72208 126756 72214
rect 126704 72150 126756 72156
rect 126624 70366 126744 70394
rect 126612 65544 126664 65550
rect 126612 65486 126664 65492
rect 126624 60110 126652 65486
rect 126716 61470 126744 70366
rect 126704 61464 126756 61470
rect 126704 61406 126756 61412
rect 126808 60178 126836 72694
rect 126900 69834 126928 75140
rect 126992 72865 127020 75140
rect 126978 72856 127034 72865
rect 126978 72791 127034 72800
rect 127084 72434 127112 75140
rect 127176 72593 127204 75140
rect 127268 72729 127296 75140
rect 127254 72720 127310 72729
rect 127254 72655 127310 72664
rect 127162 72584 127218 72593
rect 127162 72519 127218 72528
rect 127360 72457 127388 75140
rect 126992 72406 127112 72434
rect 127346 72448 127402 72457
rect 126992 71942 127020 72406
rect 127346 72383 127402 72392
rect 127452 72298 127480 75140
rect 127084 72270 127480 72298
rect 126980 71936 127032 71942
rect 126980 71878 127032 71884
rect 126888 69828 126940 69834
rect 126888 69770 126940 69776
rect 127084 66978 127112 72270
rect 127440 72208 127492 72214
rect 127440 72150 127492 72156
rect 127452 69902 127480 72150
rect 127440 69896 127492 69902
rect 127440 69838 127492 69844
rect 127072 66972 127124 66978
rect 127072 66914 127124 66920
rect 127544 65686 127572 75140
rect 127532 65680 127584 65686
rect 127532 65622 127584 65628
rect 127636 65532 127664 75140
rect 127728 72026 127756 75140
rect 127820 72214 127848 75140
rect 127912 72418 127940 75140
rect 127900 72412 127952 72418
rect 127900 72354 127952 72360
rect 127808 72208 127860 72214
rect 127808 72150 127860 72156
rect 127728 71998 127940 72026
rect 127716 71868 127768 71874
rect 127716 71810 127768 71816
rect 127452 65504 127664 65532
rect 126796 60172 126848 60178
rect 126796 60114 126848 60120
rect 126612 60104 126664 60110
rect 126612 60046 126664 60052
rect 126520 44872 126572 44878
rect 126520 44814 126572 44820
rect 127452 6254 127480 65504
rect 127728 60734 127756 71810
rect 127912 65754 127940 71998
rect 127900 65748 127952 65754
rect 127900 65690 127952 65696
rect 127808 65680 127860 65686
rect 127808 65622 127860 65628
rect 127636 60706 127756 60734
rect 127440 6248 127492 6254
rect 127440 6190 127492 6196
rect 127636 6186 127664 60706
rect 127820 57322 127848 65622
rect 127808 57316 127860 57322
rect 127808 57258 127860 57264
rect 128004 47598 128032 75140
rect 128096 71194 128124 75140
rect 128188 72350 128216 75140
rect 128176 72344 128228 72350
rect 128176 72286 128228 72292
rect 128176 71800 128228 71806
rect 128176 71742 128228 71748
rect 128084 71188 128136 71194
rect 128084 71130 128136 71136
rect 127992 47592 128044 47598
rect 127992 47534 128044 47540
rect 127624 6180 127676 6186
rect 127624 6122 127676 6128
rect 126244 3460 126296 3466
rect 126244 3402 126296 3408
rect 126980 3460 127032 3466
rect 126980 3402 127032 3408
rect 126992 480 127020 3402
rect 128188 480 128216 71742
rect 128280 65958 128308 75140
rect 128372 72865 128400 75140
rect 128358 72856 128414 72865
rect 128358 72791 128414 72800
rect 128464 72593 128492 75140
rect 128450 72584 128506 72593
rect 128450 72519 128506 72528
rect 128556 69737 128584 75140
rect 128648 72729 128676 75140
rect 128634 72720 128690 72729
rect 128634 72655 128690 72664
rect 128542 69728 128598 69737
rect 128542 69663 128598 69672
rect 128268 65952 128320 65958
rect 128268 65894 128320 65900
rect 128740 65550 128768 75140
rect 128832 68542 128860 75140
rect 128820 68536 128872 68542
rect 128820 68478 128872 68484
rect 128820 65952 128872 65958
rect 128820 65894 128872 65900
rect 128728 65544 128780 65550
rect 128728 65486 128780 65492
rect 128832 60734 128860 65894
rect 128924 65498 128952 75140
rect 129016 65958 129044 75140
rect 129108 67046 129136 75140
rect 129200 71262 129228 75140
rect 129292 73030 129320 75140
rect 129280 73024 129332 73030
rect 129280 72966 129332 72972
rect 129188 71256 129240 71262
rect 129188 71198 129240 71204
rect 129096 67040 129148 67046
rect 129096 66982 129148 66988
rect 129188 66292 129240 66298
rect 129188 66234 129240 66240
rect 129004 65952 129056 65958
rect 129004 65894 129056 65900
rect 128924 65470 129136 65498
rect 129004 65408 129056 65414
rect 129004 65350 129056 65356
rect 128832 60706 128952 60734
rect 128924 8974 128952 60706
rect 128912 8968 128964 8974
rect 128912 8910 128964 8916
rect 129016 3534 129044 65350
rect 129108 44946 129136 65470
rect 129200 65414 129228 66234
rect 129384 65822 129412 75140
rect 129372 65816 129424 65822
rect 129372 65758 129424 65764
rect 129280 65544 129332 65550
rect 129280 65486 129332 65492
rect 129188 65408 129240 65414
rect 129188 65350 129240 65356
rect 129292 47666 129320 65486
rect 129476 62966 129504 75140
rect 129568 67114 129596 75140
rect 129660 68610 129688 75140
rect 129752 73137 129780 75140
rect 129738 73128 129794 73137
rect 129738 73063 129794 73072
rect 129740 72956 129792 72962
rect 129740 72898 129792 72904
rect 129752 72078 129780 72898
rect 129844 72894 129872 75140
rect 129936 72962 129964 75140
rect 129924 72956 129976 72962
rect 129924 72898 129976 72904
rect 129832 72888 129884 72894
rect 129832 72830 129884 72836
rect 129924 72752 129976 72758
rect 129830 72720 129886 72729
rect 129924 72694 129976 72700
rect 129830 72655 129886 72664
rect 129740 72072 129792 72078
rect 129740 72014 129792 72020
rect 129844 71233 129872 72655
rect 129830 71224 129886 71233
rect 129830 71159 129886 71168
rect 129648 68604 129700 68610
rect 129648 68546 129700 68552
rect 129556 67108 129608 67114
rect 129556 67050 129608 67056
rect 129936 65890 129964 72694
rect 129924 65884 129976 65890
rect 129924 65826 129976 65832
rect 129464 62960 129516 62966
rect 129464 62902 129516 62908
rect 130028 61538 130056 75140
rect 130120 72758 130148 75140
rect 130108 72752 130160 72758
rect 130108 72694 130160 72700
rect 130108 72412 130160 72418
rect 130108 72354 130160 72360
rect 130120 68746 130148 72354
rect 130108 68740 130160 68746
rect 130108 68682 130160 68688
rect 130212 68678 130240 75140
rect 130304 72826 130332 75140
rect 130396 73098 130424 75140
rect 130384 73092 130436 73098
rect 130384 73034 130436 73040
rect 130384 72956 130436 72962
rect 130384 72898 130436 72904
rect 130292 72820 130344 72826
rect 130292 72762 130344 72768
rect 130396 70786 130424 72898
rect 130384 70780 130436 70786
rect 130384 70722 130436 70728
rect 130488 70666 130516 75140
rect 130580 72962 130608 75140
rect 130568 72956 130620 72962
rect 130568 72898 130620 72904
rect 130568 72820 130620 72826
rect 130568 72762 130620 72768
rect 130304 70638 130516 70666
rect 130200 68672 130252 68678
rect 130200 68614 130252 68620
rect 130304 67182 130332 70638
rect 130384 70508 130436 70514
rect 130384 70450 130436 70456
rect 130292 67176 130344 67182
rect 130292 67118 130344 67124
rect 130016 61532 130068 61538
rect 130016 61474 130068 61480
rect 129280 47660 129332 47666
rect 129280 47602 129332 47608
rect 129096 44940 129148 44946
rect 129096 44882 129148 44888
rect 129004 3528 129056 3534
rect 129004 3470 129056 3476
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 129384 480 129412 3470
rect 130396 2990 130424 70450
rect 130476 67652 130528 67658
rect 130476 67594 130528 67600
rect 130488 3466 130516 67594
rect 130580 64394 130608 72762
rect 130672 72418 130700 75140
rect 130660 72412 130712 72418
rect 130660 72354 130712 72360
rect 130764 70038 130792 75140
rect 130752 70032 130804 70038
rect 130752 69974 130804 69980
rect 130660 65544 130712 65550
rect 130660 65486 130712 65492
rect 130568 64388 130620 64394
rect 130568 64330 130620 64336
rect 130672 3534 130700 65486
rect 130856 60042 130884 75140
rect 130948 71330 130976 75140
rect 131040 71874 131068 75140
rect 131132 72010 131160 75140
rect 131120 72004 131172 72010
rect 131120 71946 131172 71952
rect 131028 71868 131080 71874
rect 131028 71810 131080 71816
rect 130936 71324 130988 71330
rect 130936 71266 130988 71272
rect 131224 70514 131252 75140
rect 131212 70508 131264 70514
rect 131212 70450 131264 70456
rect 131316 66298 131344 75140
rect 131408 67658 131436 75140
rect 131500 71806 131528 75140
rect 131488 71800 131540 71806
rect 131488 71742 131540 71748
rect 131396 67652 131448 67658
rect 131396 67594 131448 67600
rect 131304 66292 131356 66298
rect 131304 66234 131356 66240
rect 131592 65550 131620 75140
rect 131580 65544 131632 65550
rect 131580 65486 131632 65492
rect 131684 65226 131712 75140
rect 131776 65346 131804 75140
rect 131868 65414 131896 75140
rect 131960 65550 131988 75140
rect 131948 65544 132000 65550
rect 131948 65486 132000 65492
rect 131856 65408 131908 65414
rect 131856 65350 131908 65356
rect 131764 65340 131816 65346
rect 131764 65282 131816 65288
rect 131684 65198 131896 65226
rect 131764 65136 131816 65142
rect 131764 65078 131816 65084
rect 130844 60036 130896 60042
rect 130844 59978 130896 59984
rect 130660 3528 130712 3534
rect 130660 3470 130712 3476
rect 130476 3460 130528 3466
rect 130476 3402 130528 3408
rect 130568 3460 130620 3466
rect 130568 3402 130620 3408
rect 130384 2984 130436 2990
rect 130384 2926 130436 2932
rect 130580 480 130608 3402
rect 131776 480 131804 65078
rect 131868 60734 131896 65198
rect 131868 60706 131988 60734
rect 131960 3466 131988 60706
rect 132052 52426 132080 75140
rect 132144 65498 132172 75140
rect 132236 70394 132264 75140
rect 132328 72729 132356 75140
rect 132420 72865 132448 75140
rect 132406 72856 132462 72865
rect 132406 72791 132462 72800
rect 132314 72720 132370 72729
rect 132314 72655 132370 72664
rect 132236 70366 132448 70394
rect 132316 65544 132368 65550
rect 132144 65470 132264 65498
rect 132316 65486 132368 65492
rect 132132 65408 132184 65414
rect 132132 65350 132184 65356
rect 132040 52420 132092 52426
rect 132040 52362 132092 52368
rect 132144 42770 132172 65350
rect 132132 42764 132184 42770
rect 132132 42706 132184 42712
rect 132236 12442 132264 65470
rect 132224 12436 132276 12442
rect 132224 12378 132276 12384
rect 132328 5574 132356 65486
rect 132420 6254 132448 70366
rect 132512 65498 132540 75140
rect 132604 72350 132632 75140
rect 132592 72344 132644 72350
rect 132592 72286 132644 72292
rect 132696 72078 132724 75140
rect 132684 72072 132736 72078
rect 132684 72014 132736 72020
rect 132788 65618 132816 75140
rect 132880 66026 132908 75140
rect 132868 66020 132920 66026
rect 132868 65962 132920 65968
rect 132776 65612 132828 65618
rect 132776 65554 132828 65560
rect 132512 65470 132908 65498
rect 132592 65408 132644 65414
rect 132592 65350 132644 65356
rect 132776 65408 132828 65414
rect 132776 65350 132828 65356
rect 132604 17270 132632 65350
rect 132592 17264 132644 17270
rect 132592 17206 132644 17212
rect 132408 6248 132460 6254
rect 132408 6190 132460 6196
rect 132788 6186 132816 65350
rect 132880 60734 132908 65470
rect 132972 61962 133000 75140
rect 133064 72418 133092 75140
rect 133052 72412 133104 72418
rect 133052 72354 133104 72360
rect 133156 68474 133184 75140
rect 133144 68468 133196 68474
rect 133144 68410 133196 68416
rect 133248 62082 133276 75140
rect 133340 65634 133368 75140
rect 133432 65754 133460 75140
rect 133524 72593 133552 75140
rect 133616 72729 133644 75140
rect 133708 72865 133736 75140
rect 133694 72856 133750 72865
rect 133694 72791 133750 72800
rect 133602 72720 133658 72729
rect 133602 72655 133658 72664
rect 133510 72584 133566 72593
rect 133510 72519 133566 72528
rect 133800 72457 133828 75140
rect 133786 72448 133842 72457
rect 133604 72412 133656 72418
rect 133786 72383 133842 72392
rect 133604 72354 133656 72360
rect 133512 72344 133564 72350
rect 133512 72286 133564 72292
rect 133420 65748 133472 65754
rect 133420 65690 133472 65696
rect 133340 65606 133460 65634
rect 133432 65414 133460 65606
rect 133420 65408 133472 65414
rect 133420 65350 133472 65356
rect 133420 65272 133472 65278
rect 133420 65214 133472 65220
rect 133236 62076 133288 62082
rect 133236 62018 133288 62024
rect 132972 61934 133368 61962
rect 132880 60706 133276 60734
rect 133248 57934 133276 60706
rect 133236 57928 133288 57934
rect 133236 57870 133288 57876
rect 133340 52494 133368 61934
rect 133328 52488 133380 52494
rect 133328 52430 133380 52436
rect 133432 43450 133460 65214
rect 133420 43444 133472 43450
rect 133420 43386 133472 43392
rect 132960 42764 133012 42770
rect 132960 42706 133012 42712
rect 132776 6180 132828 6186
rect 132776 6122 132828 6128
rect 132316 5568 132368 5574
rect 132316 5510 132368 5516
rect 131948 3460 132000 3466
rect 131948 3402 132000 3408
rect 132972 480 133000 42706
rect 133524 32434 133552 72286
rect 133512 32428 133564 32434
rect 133512 32370 133564 32376
rect 133616 21418 133644 72354
rect 133892 60734 133920 75140
rect 133984 65550 134012 75140
rect 134076 73001 134104 75140
rect 134062 72992 134118 73001
rect 134062 72927 134118 72936
rect 134168 65668 134196 75140
rect 134260 65822 134288 75140
rect 134248 65816 134300 65822
rect 134248 65758 134300 65764
rect 134352 65754 134380 75140
rect 134340 65748 134392 65754
rect 134340 65690 134392 65696
rect 134168 65640 134288 65668
rect 134064 65612 134116 65618
rect 134064 65554 134116 65560
rect 133972 65544 134024 65550
rect 133972 65486 134024 65492
rect 133892 60706 134012 60734
rect 133604 21412 133656 21418
rect 133604 21354 133656 21360
rect 133984 13122 134012 60706
rect 133972 13116 134024 13122
rect 133972 13058 134024 13064
rect 133144 12436 133196 12442
rect 133144 12378 133196 12384
rect 133156 3466 133184 12378
rect 133788 5568 133840 5574
rect 133788 5510 133840 5516
rect 133144 3460 133196 3466
rect 133144 3402 133196 3408
rect 133800 2802 133828 5510
rect 134076 3398 134104 65554
rect 134260 60734 134288 65640
rect 134444 65618 134472 75140
rect 134536 72162 134564 75140
rect 134628 72758 134656 75140
rect 134616 72752 134668 72758
rect 134616 72694 134668 72700
rect 134536 72134 134656 72162
rect 134524 72072 134576 72078
rect 134524 72014 134576 72020
rect 134432 65612 134484 65618
rect 134432 65554 134484 65560
rect 134260 60706 134472 60734
rect 134444 40730 134472 60706
rect 134432 40724 134484 40730
rect 134432 40666 134484 40672
rect 134536 4826 134564 72014
rect 134628 68882 134656 72134
rect 134720 70174 134748 75140
rect 134812 72457 134840 75140
rect 134904 72729 134932 75140
rect 134996 74361 135024 75140
rect 134982 74352 135038 74361
rect 134982 74287 135038 74296
rect 135088 72865 135116 75140
rect 135074 72856 135130 72865
rect 135074 72791 135130 72800
rect 135076 72752 135128 72758
rect 134890 72720 134946 72729
rect 135076 72694 135128 72700
rect 134890 72655 134946 72664
rect 134798 72448 134854 72457
rect 134798 72383 134854 72392
rect 134708 70168 134760 70174
rect 134708 70110 134760 70116
rect 134616 68876 134668 68882
rect 134616 68818 134668 68824
rect 134616 66020 134668 66026
rect 134616 65962 134668 65968
rect 134524 4820 134576 4826
rect 134524 4762 134576 4768
rect 134628 3738 134656 65962
rect 135088 65822 135116 72694
rect 135180 72593 135208 75140
rect 135166 72584 135222 72593
rect 135166 72519 135222 72528
rect 134892 65816 134944 65822
rect 134892 65758 134944 65764
rect 135076 65816 135128 65822
rect 135076 65758 135128 65764
rect 134800 65748 134852 65754
rect 134800 65690 134852 65696
rect 134708 52420 134760 52426
rect 134708 52362 134760 52368
rect 134616 3732 134668 3738
rect 134616 3674 134668 3680
rect 134720 3534 134748 52362
rect 134812 36650 134840 65690
rect 134800 36644 134852 36650
rect 134800 36586 134852 36592
rect 134904 31074 134932 65758
rect 134984 65544 135036 65550
rect 134984 65486 135036 65492
rect 134892 31068 134944 31074
rect 134892 31010 134944 31016
rect 134996 29782 135024 65486
rect 135272 58954 135300 75140
rect 135364 65414 135392 75140
rect 135456 74905 135484 75140
rect 135442 74896 135498 74905
rect 135442 74831 135498 74840
rect 135444 74792 135496 74798
rect 135444 74734 135496 74740
rect 135456 74594 135484 74734
rect 135444 74588 135496 74594
rect 135444 74530 135496 74536
rect 135444 72140 135496 72146
rect 135444 72082 135496 72088
rect 135456 68814 135484 72082
rect 135444 68808 135496 68814
rect 135444 68750 135496 68756
rect 135352 65408 135404 65414
rect 135352 65350 135404 65356
rect 135548 60734 135576 75140
rect 135640 72146 135668 75140
rect 135628 72140 135680 72146
rect 135628 72082 135680 72088
rect 135628 65612 135680 65618
rect 135628 65554 135680 65560
rect 135456 60706 135576 60734
rect 135260 58948 135312 58954
rect 135260 58890 135312 58896
rect 135456 47870 135484 60706
rect 135444 47864 135496 47870
rect 135444 47806 135496 47812
rect 135640 46306 135668 65554
rect 135732 64326 135760 75140
rect 135720 64320 135772 64326
rect 135720 64262 135772 64268
rect 135628 46300 135680 46306
rect 135628 46242 135680 46248
rect 135824 39574 135852 75140
rect 135916 72350 135944 75140
rect 135904 72344 135956 72350
rect 135904 72286 135956 72292
rect 135904 68468 135956 68474
rect 135904 68410 135956 68416
rect 135812 39568 135864 39574
rect 135812 39510 135864 39516
rect 134984 29776 135036 29782
rect 134984 29718 135036 29724
rect 135916 3670 135944 68410
rect 136008 65498 136036 75140
rect 136100 70854 136128 75140
rect 136088 70848 136140 70854
rect 136088 70790 136140 70796
rect 136192 65618 136220 75140
rect 136284 72457 136312 75140
rect 136376 72729 136404 75140
rect 136468 72865 136496 75140
rect 136454 72856 136510 72865
rect 136454 72791 136510 72800
rect 136362 72720 136418 72729
rect 136362 72655 136418 72664
rect 136560 72593 136588 75140
rect 136652 73030 136680 75140
rect 136640 73024 136692 73030
rect 136640 72966 136692 72972
rect 136546 72584 136602 72593
rect 136546 72519 136602 72528
rect 136270 72448 136326 72457
rect 136270 72383 136326 72392
rect 136272 72344 136324 72350
rect 136272 72286 136324 72292
rect 136180 65612 136232 65618
rect 136180 65554 136232 65560
rect 136008 65470 136220 65498
rect 136088 65408 136140 65414
rect 136088 65350 136140 65356
rect 135996 62076 136048 62082
rect 135996 62018 136048 62024
rect 135904 3664 135956 3670
rect 135904 3606 135956 3612
rect 136008 3602 136036 62018
rect 136100 56030 136128 65350
rect 136088 56024 136140 56030
rect 136088 55966 136140 55972
rect 136192 53514 136220 65470
rect 136180 53508 136232 53514
rect 136180 53450 136232 53456
rect 136180 52488 136232 52494
rect 136180 52430 136232 52436
rect 136192 3806 136220 52430
rect 136284 49094 136312 72286
rect 136744 62966 136772 75140
rect 136836 72321 136864 75140
rect 136822 72312 136878 72321
rect 136822 72247 136878 72256
rect 136824 65680 136876 65686
rect 136824 65622 136876 65628
rect 136732 62960 136784 62966
rect 136732 62902 136784 62908
rect 136364 57928 136416 57934
rect 136364 57870 136416 57876
rect 136272 49088 136324 49094
rect 136272 49030 136324 49036
rect 136270 48240 136326 48249
rect 136270 48175 136326 48184
rect 136180 3800 136232 3806
rect 136180 3742 136232 3748
rect 135996 3596 136048 3602
rect 135996 3538 136048 3544
rect 136284 3534 136312 48175
rect 134708 3528 134760 3534
rect 134708 3470 134760 3476
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 136272 3528 136324 3534
rect 136272 3470 136324 3476
rect 134064 3392 134116 3398
rect 134064 3334 134116 3340
rect 133800 2774 133920 2802
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 2774
rect 135272 480 135300 3470
rect 136376 2990 136404 57870
rect 136836 6118 136864 65622
rect 136928 65550 136956 75140
rect 136916 65544 136968 65550
rect 136916 65486 136968 65492
rect 136824 6112 136876 6118
rect 136824 6054 136876 6060
rect 137020 5166 137048 75140
rect 137112 66774 137140 75140
rect 137100 66768 137152 66774
rect 137100 66710 137152 66716
rect 137100 65748 137152 65754
rect 137100 65690 137152 65696
rect 137112 60734 137140 65690
rect 137204 65498 137232 75140
rect 137296 65618 137324 75140
rect 137284 65612 137336 65618
rect 137284 65554 137336 65560
rect 137204 65470 137324 65498
rect 137112 60706 137232 60734
rect 137204 60246 137232 60706
rect 137192 60240 137244 60246
rect 137192 60182 137244 60188
rect 137296 53446 137324 65470
rect 137284 53440 137336 53446
rect 137284 53382 137336 53388
rect 137388 50658 137416 75140
rect 137480 65686 137508 75140
rect 137468 65680 137520 65686
rect 137468 65622 137520 65628
rect 137468 65544 137520 65550
rect 137468 65486 137520 65492
rect 137376 50652 137428 50658
rect 137376 50594 137428 50600
rect 137480 43654 137508 65486
rect 137468 43648 137520 43654
rect 137468 43590 137520 43596
rect 137572 38146 137600 75140
rect 137664 65754 137692 75140
rect 137756 71505 137784 75140
rect 137848 72729 137876 75140
rect 137940 72865 137968 75140
rect 137926 72856 137982 72865
rect 137926 72791 137982 72800
rect 137834 72720 137890 72729
rect 137834 72655 137890 72664
rect 137742 71496 137798 71505
rect 137742 71431 137798 71440
rect 137744 66768 137796 66774
rect 137744 66710 137796 66716
rect 137652 65748 137704 65754
rect 137652 65690 137704 65696
rect 137652 65612 137704 65618
rect 137652 65554 137704 65560
rect 137560 38140 137612 38146
rect 137560 38082 137612 38088
rect 137664 18834 137692 65554
rect 137756 63102 137784 66710
rect 138032 65142 138060 75140
rect 138124 72146 138152 75140
rect 138112 72140 138164 72146
rect 138112 72082 138164 72088
rect 138216 71913 138244 75140
rect 138202 71904 138258 71913
rect 138202 71839 138258 71848
rect 138308 70394 138336 75140
rect 138216 70366 138336 70394
rect 138020 65136 138072 65142
rect 138020 65078 138072 65084
rect 138216 65006 138244 70366
rect 138400 65686 138428 75140
rect 138492 72185 138520 75140
rect 138478 72176 138534 72185
rect 138478 72111 138534 72120
rect 138584 65686 138612 75140
rect 138388 65680 138440 65686
rect 138388 65622 138440 65628
rect 138572 65680 138624 65686
rect 138572 65622 138624 65628
rect 138676 65498 138704 75140
rect 138768 65958 138796 75140
rect 138756 65952 138808 65958
rect 138756 65894 138808 65900
rect 138308 65470 138704 65498
rect 138204 65000 138256 65006
rect 138204 64942 138256 64948
rect 137744 63096 137796 63102
rect 137744 63038 137796 63044
rect 137744 62960 137796 62966
rect 137744 62902 137796 62908
rect 137652 18828 137704 18834
rect 137652 18770 137704 18776
rect 137652 6248 137704 6254
rect 137652 6190 137704 6196
rect 137008 5160 137060 5166
rect 137008 5102 137060 5108
rect 136456 3460 136508 3466
rect 136456 3402 136508 3408
rect 136364 2984 136416 2990
rect 136364 2926 136416 2932
rect 136468 480 136496 3402
rect 137664 480 137692 6190
rect 137756 6050 137784 62902
rect 138308 17542 138336 65470
rect 138860 65362 138888 75140
rect 138952 65550 138980 75140
rect 138940 65544 138992 65550
rect 138940 65486 138992 65492
rect 138492 65334 138888 65362
rect 138940 65408 138992 65414
rect 138940 65350 138992 65356
rect 138296 17536 138348 17542
rect 138296 17478 138348 17484
rect 138492 16182 138520 65334
rect 138664 65272 138716 65278
rect 138664 65214 138716 65220
rect 138676 57458 138704 65214
rect 138756 65204 138808 65210
rect 138756 65146 138808 65152
rect 138664 57452 138716 57458
rect 138664 57394 138716 57400
rect 138768 54806 138796 65146
rect 138848 65136 138900 65142
rect 138848 65078 138900 65084
rect 138952 65090 138980 65350
rect 139044 65278 139072 75140
rect 139136 73545 139164 75140
rect 139122 73536 139178 73545
rect 139122 73471 139178 73480
rect 139228 73409 139256 75140
rect 139214 73400 139270 73409
rect 139214 73335 139270 73344
rect 139320 73137 139348 75140
rect 139306 73128 139362 73137
rect 139306 73063 139362 73072
rect 139308 72140 139360 72146
rect 139308 72082 139360 72088
rect 139320 68746 139348 72082
rect 139308 68740 139360 68746
rect 139308 68682 139360 68688
rect 139216 65952 139268 65958
rect 139216 65894 139268 65900
rect 139124 65544 139176 65550
rect 139124 65486 139176 65492
rect 139032 65272 139084 65278
rect 139032 65214 139084 65220
rect 138756 54800 138808 54806
rect 138756 54742 138808 54748
rect 138860 42294 138888 65078
rect 138952 65062 139072 65090
rect 138940 65000 138992 65006
rect 138940 64942 138992 64948
rect 138848 42288 138900 42294
rect 138848 42230 138900 42236
rect 138952 40934 138980 64942
rect 138940 40928 138992 40934
rect 138940 40870 138992 40876
rect 139044 32706 139072 65062
rect 139032 32700 139084 32706
rect 139032 32642 139084 32648
rect 139136 28626 139164 65486
rect 139228 61538 139256 65894
rect 139412 65686 139440 75140
rect 139400 65680 139452 65686
rect 139400 65622 139452 65628
rect 139504 65550 139532 75140
rect 139596 74225 139624 75140
rect 139582 74216 139638 74225
rect 139582 74151 139638 74160
rect 139584 73976 139636 73982
rect 139584 73918 139636 73924
rect 139596 72457 139624 73918
rect 139582 72448 139638 72457
rect 139582 72383 139638 72392
rect 139688 70394 139716 75140
rect 139596 70366 139716 70394
rect 139492 65544 139544 65550
rect 139492 65486 139544 65492
rect 139596 65278 139624 70366
rect 139780 65754 139808 75140
rect 139872 73273 139900 75140
rect 139858 73264 139914 73273
rect 139858 73199 139914 73208
rect 139860 73024 139912 73030
rect 139860 72966 139912 72972
rect 139872 70990 139900 72966
rect 139860 70984 139912 70990
rect 139860 70926 139912 70932
rect 139964 65890 139992 75140
rect 139952 65884 140004 65890
rect 139952 65826 140004 65832
rect 139768 65748 139820 65754
rect 139768 65690 139820 65696
rect 140056 65600 140084 75140
rect 139688 65572 140084 65600
rect 139584 65272 139636 65278
rect 139584 65214 139636 65220
rect 139216 61532 139268 61538
rect 139216 61474 139268 61480
rect 139124 28620 139176 28626
rect 139124 28562 139176 28568
rect 139688 18766 139716 65572
rect 139860 65476 139912 65482
rect 139860 65418 139912 65424
rect 139676 18760 139728 18766
rect 139676 18702 139728 18708
rect 138480 16176 138532 16182
rect 138480 16118 138532 16124
rect 139872 13394 139900 65418
rect 140148 60178 140176 75140
rect 140240 65482 140268 75140
rect 140332 68678 140360 75140
rect 140424 73409 140452 75140
rect 140516 73545 140544 75140
rect 140502 73536 140558 73545
rect 140502 73471 140558 73480
rect 140608 73409 140636 75140
rect 140700 73681 140728 75140
rect 140792 73846 140820 75140
rect 140780 73840 140832 73846
rect 140780 73782 140832 73788
rect 140686 73672 140742 73681
rect 140686 73607 140742 73616
rect 140780 73636 140832 73642
rect 140780 73578 140832 73584
rect 140410 73400 140466 73409
rect 140410 73335 140466 73344
rect 140594 73400 140650 73409
rect 140594 73335 140650 73344
rect 140792 71670 140820 73578
rect 140780 71664 140832 71670
rect 140780 71606 140832 71612
rect 140320 68672 140372 68678
rect 140320 68614 140372 68620
rect 140412 65884 140464 65890
rect 140412 65826 140464 65832
rect 140320 65748 140372 65754
rect 140320 65690 140372 65696
rect 140228 65476 140280 65482
rect 140228 65418 140280 65424
rect 140332 65362 140360 65690
rect 140240 65334 140360 65362
rect 140136 60172 140188 60178
rect 140136 60114 140188 60120
rect 140240 46238 140268 65334
rect 140320 65272 140372 65278
rect 140320 65214 140372 65220
rect 140228 46232 140280 46238
rect 140228 46174 140280 46180
rect 140332 31346 140360 65214
rect 140320 31340 140372 31346
rect 140320 31282 140372 31288
rect 140424 24478 140452 65826
rect 140884 65550 140912 75140
rect 140976 73710 141004 75140
rect 140964 73704 141016 73710
rect 140964 73646 141016 73652
rect 141068 73642 141096 75140
rect 141056 73636 141108 73642
rect 141056 73578 141108 73584
rect 141160 73522 141188 75140
rect 140964 73500 141016 73506
rect 140964 73442 141016 73448
rect 141068 73494 141188 73522
rect 141252 73506 141280 75140
rect 141240 73500 141292 73506
rect 140976 71602 141004 73442
rect 140964 71596 141016 71602
rect 140964 71538 141016 71544
rect 141068 68134 141096 73494
rect 141240 73442 141292 73448
rect 141148 73432 141200 73438
rect 141148 73374 141200 73380
rect 141056 68128 141108 68134
rect 141056 68070 141108 68076
rect 140504 65544 140556 65550
rect 140504 65486 140556 65492
rect 140872 65544 140924 65550
rect 140872 65486 140924 65492
rect 140412 24472 140464 24478
rect 140412 24414 140464 24420
rect 140516 21690 140544 65486
rect 140504 21684 140556 21690
rect 140504 21626 140556 21632
rect 140042 17232 140098 17241
rect 140042 17167 140098 17176
rect 139860 13388 139912 13394
rect 139860 13330 139912 13336
rect 137744 6044 137796 6050
rect 137744 5986 137796 5992
rect 138846 3360 138902 3369
rect 138846 3295 138902 3304
rect 138860 480 138888 3295
rect 140056 480 140084 17167
rect 141160 4146 141188 73374
rect 141240 73364 141292 73370
rect 141240 73306 141292 73312
rect 141252 71774 141280 73306
rect 141344 71890 141372 75140
rect 141436 73982 141464 75140
rect 141424 73976 141476 73982
rect 141424 73918 141476 73924
rect 141424 73840 141476 73846
rect 141424 73782 141476 73788
rect 141436 73166 141464 73782
rect 141528 73438 141556 75140
rect 141516 73432 141568 73438
rect 141516 73374 141568 73380
rect 141424 73160 141476 73166
rect 141424 73102 141476 73108
rect 141620 72690 141648 75140
rect 141712 73642 141740 75140
rect 141700 73636 141752 73642
rect 141700 73578 141752 73584
rect 141804 73522 141832 75140
rect 141712 73494 141832 73522
rect 141608 72684 141660 72690
rect 141608 72626 141660 72632
rect 141344 71862 141648 71890
rect 141252 71746 141372 71774
rect 141344 70394 141372 71746
rect 141344 70366 141464 70394
rect 141240 67040 141292 67046
rect 141240 66982 141292 66988
rect 141148 4140 141200 4146
rect 141148 4082 141200 4088
rect 141252 4078 141280 66982
rect 141436 36718 141464 70366
rect 141516 68128 141568 68134
rect 141516 68070 141568 68076
rect 141424 36712 141476 36718
rect 141424 36654 141476 36660
rect 141528 6798 141556 68070
rect 141516 6792 141568 6798
rect 141516 6734 141568 6740
rect 141620 6730 141648 71862
rect 141712 67046 141740 73494
rect 141792 72684 141844 72690
rect 141792 72626 141844 72632
rect 141700 67040 141752 67046
rect 141700 66982 141752 66988
rect 141700 66904 141752 66910
rect 141700 66846 141752 66852
rect 141608 6724 141660 6730
rect 141608 6666 141660 6672
rect 141712 6594 141740 66846
rect 141804 66756 141832 72626
rect 141896 66910 141924 75140
rect 141988 69737 142016 75140
rect 142080 73545 142108 75140
rect 142066 73536 142122 73545
rect 142066 73471 142122 73480
rect 142068 73432 142120 73438
rect 142068 73374 142120 73380
rect 142080 72321 142108 73374
rect 142066 72312 142122 72321
rect 142066 72247 142122 72256
rect 141974 69728 142030 69737
rect 141974 69663 142030 69672
rect 141884 66904 141936 66910
rect 141884 66846 141936 66852
rect 141804 66728 141924 66756
rect 141792 65544 141844 65550
rect 141792 65486 141844 65492
rect 141804 6866 141832 65486
rect 141792 6860 141844 6866
rect 141792 6802 141844 6808
rect 141896 6662 141924 66728
rect 142172 7818 142200 75140
rect 142264 65618 142292 75140
rect 142356 74089 142384 75140
rect 142342 74080 142398 74089
rect 142342 74015 142398 74024
rect 142344 73160 142396 73166
rect 142344 73102 142396 73108
rect 142356 71058 142384 73102
rect 142344 71052 142396 71058
rect 142344 70994 142396 71000
rect 142252 65612 142304 65618
rect 142252 65554 142304 65560
rect 142448 65550 142476 75140
rect 142436 65544 142488 65550
rect 142436 65486 142488 65492
rect 142540 65278 142568 75140
rect 142528 65272 142580 65278
rect 142528 65214 142580 65220
rect 142632 60734 142660 75140
rect 142724 65958 142752 75140
rect 142816 67522 142844 75140
rect 142804 67516 142856 67522
rect 142804 67458 142856 67464
rect 142712 65952 142764 65958
rect 142712 65894 142764 65900
rect 142908 65532 142936 75140
rect 143000 70394 143028 75140
rect 143092 73166 143120 75140
rect 143080 73160 143132 73166
rect 143080 73102 143132 73108
rect 143184 72729 143212 75140
rect 143276 72865 143304 75140
rect 143368 73001 143396 75140
rect 143354 72992 143410 73001
rect 143354 72927 143410 72936
rect 143262 72856 143318 72865
rect 143262 72791 143318 72800
rect 143170 72720 143226 72729
rect 143170 72655 143226 72664
rect 143460 72593 143488 75140
rect 143446 72584 143502 72593
rect 143446 72519 143502 72528
rect 143552 71534 143580 75140
rect 143540 71528 143592 71534
rect 143540 71470 143592 71476
rect 143000 70366 143396 70394
rect 143080 67516 143132 67522
rect 143080 67458 143132 67464
rect 142988 65952 143040 65958
rect 142988 65894 143040 65900
rect 142724 65504 142936 65532
rect 142724 65260 142752 65504
rect 142896 65272 142948 65278
rect 142724 65232 142844 65260
rect 142632 60706 142752 60734
rect 142724 57390 142752 60706
rect 142712 57384 142764 57390
rect 142712 57326 142764 57332
rect 142816 54738 142844 65232
rect 142896 65214 142948 65220
rect 142804 54732 142856 54738
rect 142804 54674 142856 54680
rect 142908 40866 142936 65214
rect 142896 40860 142948 40866
rect 142896 40802 142948 40808
rect 143000 35426 143028 65894
rect 142988 35420 143040 35426
rect 142988 35362 143040 35368
rect 143092 33930 143120 67458
rect 143264 65612 143316 65618
rect 143264 65554 143316 65560
rect 143172 65544 143224 65550
rect 143172 65486 143224 65492
rect 143080 33924 143132 33930
rect 143080 33866 143132 33872
rect 142436 32428 142488 32434
rect 142436 32370 142488 32376
rect 142160 7812 142212 7818
rect 142160 7754 142212 7760
rect 141884 6656 141936 6662
rect 141884 6598 141936 6604
rect 141700 6588 141752 6594
rect 141700 6530 141752 6536
rect 141240 4072 141292 4078
rect 141240 4014 141292 4020
rect 141240 2984 141292 2990
rect 141240 2926 141292 2932
rect 141252 480 141280 2926
rect 142448 480 142476 32370
rect 143184 28558 143212 65486
rect 143172 28552 143224 28558
rect 143172 28494 143224 28500
rect 143276 20262 143304 65554
rect 143264 20256 143316 20262
rect 143264 20198 143316 20204
rect 143368 14754 143396 70366
rect 143644 65618 143672 75140
rect 143736 74934 143764 75140
rect 143724 74928 143776 74934
rect 143724 74870 143776 74876
rect 143724 74792 143776 74798
rect 143724 74734 143776 74740
rect 143736 72321 143764 74734
rect 143722 72312 143778 72321
rect 143722 72247 143778 72256
rect 143632 65612 143684 65618
rect 143632 65554 143684 65560
rect 143828 39506 143856 75140
rect 143920 65414 143948 75140
rect 144012 71466 144040 75140
rect 144000 71460 144052 71466
rect 144000 71402 144052 71408
rect 144000 65680 144052 65686
rect 144000 65622 144052 65628
rect 143908 65408 143960 65414
rect 143908 65350 143960 65356
rect 143816 39500 143868 39506
rect 143816 39442 143868 39448
rect 143356 14748 143408 14754
rect 143356 14690 143408 14696
rect 143540 4820 143592 4826
rect 143540 4762 143592 4768
rect 143552 480 143580 4762
rect 144012 3942 144040 65622
rect 144104 65550 144132 75140
rect 144092 65544 144144 65550
rect 144092 65486 144144 65492
rect 144196 47802 144224 75140
rect 144288 65686 144316 75140
rect 144276 65680 144328 65686
rect 144276 65622 144328 65628
rect 144380 65532 144408 75140
rect 144288 65504 144408 65532
rect 144184 47796 144236 47802
rect 144184 47738 144236 47744
rect 144288 32638 144316 65504
rect 144368 65408 144420 65414
rect 144368 65350 144420 65356
rect 144276 32632 144328 32638
rect 144276 32574 144328 32580
rect 144380 22914 144408 65350
rect 144368 22908 144420 22914
rect 144368 22850 144420 22856
rect 144472 20126 144500 75140
rect 144564 72457 144592 75140
rect 144656 72593 144684 75140
rect 144748 72729 144776 75140
rect 144840 72865 144868 75140
rect 144826 72856 144882 72865
rect 144826 72791 144882 72800
rect 144734 72720 144790 72729
rect 144734 72655 144790 72664
rect 144642 72584 144698 72593
rect 144642 72519 144698 72528
rect 144826 72584 144882 72593
rect 144826 72519 144882 72528
rect 144550 72448 144606 72457
rect 144550 72383 144606 72392
rect 144840 72185 144868 72519
rect 144826 72176 144882 72185
rect 144826 72111 144882 72120
rect 144932 65618 144960 75140
rect 144552 65612 144604 65618
rect 144552 65554 144604 65560
rect 144920 65612 144972 65618
rect 144920 65554 144972 65560
rect 144564 20194 144592 65554
rect 144644 65544 144696 65550
rect 144644 65486 144696 65492
rect 144552 20188 144604 20194
rect 144552 20130 144604 20136
rect 144460 20120 144512 20126
rect 144460 20062 144512 20068
rect 144656 14686 144684 65486
rect 144736 43444 144788 43450
rect 144736 43386 144788 43392
rect 144644 14680 144696 14686
rect 144644 14622 144696 14628
rect 144000 3936 144052 3942
rect 144000 3878 144052 3884
rect 144748 480 144776 43386
rect 145024 6526 145052 75140
rect 145116 72894 145144 75140
rect 145104 72888 145156 72894
rect 145104 72830 145156 72836
rect 145104 72752 145156 72758
rect 145104 72694 145156 72700
rect 145116 9246 145144 72694
rect 145208 65550 145236 75140
rect 145300 70394 145328 75140
rect 145392 73001 145420 75140
rect 145378 72992 145434 73001
rect 145378 72927 145434 72936
rect 145484 71398 145512 75140
rect 145472 71392 145524 71398
rect 145472 71334 145524 71340
rect 145576 70922 145604 75140
rect 145564 70916 145616 70922
rect 145564 70858 145616 70864
rect 145300 70366 145420 70394
rect 145196 65544 145248 65550
rect 145196 65486 145248 65492
rect 145104 9240 145156 9246
rect 145104 9182 145156 9188
rect 145012 6520 145064 6526
rect 145012 6462 145064 6468
rect 145392 6458 145420 70366
rect 145564 66904 145616 66910
rect 145564 66846 145616 66852
rect 145576 57322 145604 66846
rect 145564 57316 145616 57322
rect 145564 57258 145616 57264
rect 145668 50590 145696 75140
rect 145760 70242 145788 75140
rect 145852 72758 145880 75140
rect 145840 72752 145892 72758
rect 145840 72694 145892 72700
rect 145840 70916 145892 70922
rect 145840 70858 145892 70864
rect 145748 70236 145800 70242
rect 145748 70178 145800 70184
rect 145852 66756 145880 70858
rect 145944 66910 145972 75140
rect 146036 71806 146064 75140
rect 146128 72729 146156 75140
rect 146220 72865 146248 75140
rect 146206 72856 146262 72865
rect 146206 72791 146262 72800
rect 146114 72720 146170 72729
rect 146114 72655 146170 72664
rect 146024 71800 146076 71806
rect 146024 71742 146076 71748
rect 145932 66904 145984 66910
rect 145932 66846 145984 66852
rect 145852 66728 145972 66756
rect 145748 65612 145800 65618
rect 145748 65554 145800 65560
rect 145656 50584 145708 50590
rect 145656 50526 145708 50532
rect 145760 38078 145788 65554
rect 145840 65544 145892 65550
rect 145840 65486 145892 65492
rect 145748 38072 145800 38078
rect 145748 38014 145800 38020
rect 145852 25770 145880 65486
rect 145840 25764 145892 25770
rect 145840 25706 145892 25712
rect 145944 9314 145972 66728
rect 146312 65278 146340 75140
rect 146300 65272 146352 65278
rect 146300 65214 146352 65220
rect 146404 63782 146432 75140
rect 146496 74934 146524 75140
rect 146484 74928 146536 74934
rect 146484 74870 146536 74876
rect 146392 63776 146444 63782
rect 146392 63718 146444 63724
rect 146588 60734 146616 75140
rect 146680 65414 146708 75140
rect 146668 65408 146720 65414
rect 146668 65350 146720 65356
rect 146496 60706 146616 60734
rect 146772 60734 146800 75140
rect 146864 65346 146892 75140
rect 146956 67114 146984 75140
rect 146944 67108 146996 67114
rect 146944 67050 146996 67056
rect 146852 65340 146904 65346
rect 146852 65282 146904 65288
rect 147048 63866 147076 75140
rect 147140 65532 147168 75140
rect 147232 70394 147260 75140
rect 147324 72729 147352 75140
rect 147310 72720 147366 72729
rect 147310 72655 147366 72664
rect 147416 72185 147444 75140
rect 147402 72176 147458 72185
rect 147402 72111 147458 72120
rect 147508 71505 147536 75140
rect 147494 71496 147550 71505
rect 147494 71431 147550 71440
rect 147600 71369 147628 75140
rect 147586 71360 147642 71369
rect 147586 71295 147642 71304
rect 147232 70366 147536 70394
rect 147140 65504 147444 65532
rect 147220 65408 147272 65414
rect 147220 65350 147272 65356
rect 147128 65272 147180 65278
rect 147128 65214 147180 65220
rect 146956 63838 147076 63866
rect 146772 60706 146892 60734
rect 145932 9308 145984 9314
rect 145932 9250 145984 9256
rect 145380 6452 145432 6458
rect 145380 6394 145432 6400
rect 146496 5098 146524 60706
rect 146864 54670 146892 60706
rect 146852 54664 146904 54670
rect 146852 54606 146904 54612
rect 146956 51950 146984 63838
rect 147036 63776 147088 63782
rect 147036 63718 147088 63724
rect 146944 51944 146996 51950
rect 146944 51886 146996 51892
rect 147048 35358 147076 63718
rect 147036 35352 147088 35358
rect 147036 35294 147088 35300
rect 147140 24410 147168 65214
rect 147128 24404 147180 24410
rect 147128 24346 147180 24352
rect 147232 16114 147260 65350
rect 147312 65340 147364 65346
rect 147312 65282 147364 65288
rect 147220 16108 147272 16114
rect 147220 16050 147272 16056
rect 147324 13326 147352 65282
rect 147312 13320 147364 13326
rect 147312 13262 147364 13268
rect 147416 10538 147444 65504
rect 147404 10532 147456 10538
rect 147404 10474 147456 10480
rect 146484 5092 146536 5098
rect 146484 5034 146536 5040
rect 147508 5030 147536 70366
rect 147692 65550 147720 75140
rect 147784 73098 147812 75140
rect 147772 73092 147824 73098
rect 147772 73034 147824 73040
rect 147770 72992 147826 73001
rect 147770 72927 147826 72936
rect 147784 72185 147812 72927
rect 147770 72176 147826 72185
rect 147770 72111 147826 72120
rect 147680 65544 147732 65550
rect 147680 65486 147732 65492
rect 147876 65278 147904 75140
rect 147864 65272 147916 65278
rect 147864 65214 147916 65220
rect 147968 7750 147996 75140
rect 148060 65618 148088 75140
rect 148152 70394 148180 75140
rect 148244 74458 148272 75140
rect 148232 74452 148284 74458
rect 148232 74394 148284 74400
rect 148232 74316 148284 74322
rect 148232 74258 148284 74264
rect 148244 74118 148272 74258
rect 148232 74112 148284 74118
rect 148232 74054 148284 74060
rect 148232 73092 148284 73098
rect 148232 73034 148284 73040
rect 148244 72418 148272 73034
rect 148232 72412 148284 72418
rect 148232 72354 148284 72360
rect 148152 70366 148272 70394
rect 148048 65612 148100 65618
rect 148048 65554 148100 65560
rect 148140 65544 148192 65550
rect 148140 65486 148192 65492
rect 148152 14618 148180 65486
rect 148244 65362 148272 70366
rect 148336 65550 148364 75140
rect 148324 65544 148376 65550
rect 148324 65486 148376 65492
rect 148428 65498 148456 75140
rect 148520 69630 148548 75140
rect 148612 72570 148640 75140
rect 148704 73137 148732 75140
rect 148690 73128 148746 73137
rect 148690 73063 148746 73072
rect 148796 72729 148824 75140
rect 148888 72865 148916 75140
rect 148874 72856 148930 72865
rect 148874 72791 148930 72800
rect 148782 72720 148838 72729
rect 148782 72655 148838 72664
rect 148980 72593 149008 75140
rect 148966 72584 149022 72593
rect 148612 72542 148916 72570
rect 148600 72412 148652 72418
rect 148600 72354 148652 72360
rect 148508 69624 148560 69630
rect 148508 69566 148560 69572
rect 148428 65470 148548 65498
rect 148244 65334 148456 65362
rect 148324 65272 148376 65278
rect 148324 65214 148376 65220
rect 148336 60110 148364 65214
rect 148324 60104 148376 60110
rect 148324 60046 148376 60052
rect 148428 53378 148456 65334
rect 148416 53372 148468 53378
rect 148416 53314 148468 53320
rect 148520 49026 148548 65470
rect 148508 49020 148560 49026
rect 148508 48962 148560 48968
rect 148612 32570 148640 72354
rect 148888 67046 148916 72542
rect 148966 72519 149022 72528
rect 149072 71874 149100 75140
rect 149164 72214 149192 75140
rect 149152 72208 149204 72214
rect 149152 72150 149204 72156
rect 149060 71868 149112 71874
rect 149060 71810 149112 71816
rect 149256 70394 149284 75140
rect 149072 70366 149284 70394
rect 148876 67040 148928 67046
rect 148876 66982 148928 66988
rect 148784 65612 148836 65618
rect 148784 65554 148836 65560
rect 148692 65544 148744 65550
rect 148692 65486 148744 65492
rect 148600 32564 148652 32570
rect 148600 32506 148652 32512
rect 148704 21554 148732 65486
rect 148796 21622 148824 65554
rect 149072 62966 149100 70366
rect 149348 65686 149376 75140
rect 149336 65680 149388 65686
rect 149336 65622 149388 65628
rect 149440 65498 149468 75140
rect 149164 65470 149468 65498
rect 149060 62960 149112 62966
rect 149060 62902 149112 62908
rect 148784 21616 148836 21622
rect 148784 21558 148836 21564
rect 148692 21548 148744 21554
rect 148692 21490 148744 21496
rect 149164 21486 149192 65470
rect 149428 65408 149480 65414
rect 149242 65376 149298 65385
rect 149428 65350 149480 65356
rect 149242 65311 149298 65320
rect 149152 21480 149204 21486
rect 149152 21422 149204 21428
rect 149256 21418 149284 65311
rect 148324 21412 148376 21418
rect 148324 21354 148376 21360
rect 149244 21412 149296 21418
rect 149244 21354 149296 21360
rect 148140 14612 148192 14618
rect 148140 14554 148192 14560
rect 147956 7744 148008 7750
rect 147956 7686 148008 7692
rect 147496 5024 147548 5030
rect 147496 4966 147548 4972
rect 147128 3800 147180 3806
rect 147128 3742 147180 3748
rect 145932 3732 145984 3738
rect 145932 3674 145984 3680
rect 145944 480 145972 3674
rect 147140 480 147168 3742
rect 148336 480 148364 21354
rect 149440 9178 149468 65350
rect 149532 60734 149560 75140
rect 149624 65550 149652 75140
rect 149716 72350 149744 75140
rect 149704 72344 149756 72350
rect 149704 72286 149756 72292
rect 149704 71800 149756 71806
rect 149704 71742 149756 71748
rect 149612 65544 149664 65550
rect 149612 65486 149664 65492
rect 149532 60706 149652 60734
rect 149624 55962 149652 60706
rect 149612 55956 149664 55962
rect 149612 55898 149664 55904
rect 149716 27130 149744 71742
rect 149808 65498 149836 75140
rect 149900 65618 149928 75140
rect 149992 65657 150020 75140
rect 149978 65648 150034 65657
rect 149888 65612 149940 65618
rect 149978 65583 150034 65592
rect 149888 65554 149940 65560
rect 149980 65544 150032 65550
rect 149808 65470 149928 65498
rect 149980 65486 150032 65492
rect 149796 61124 149848 61130
rect 149796 61066 149848 61072
rect 149808 50522 149836 61066
rect 149796 50516 149848 50522
rect 149796 50458 149848 50464
rect 149900 47734 149928 65470
rect 149888 47728 149940 47734
rect 149888 47670 149940 47676
rect 149992 42226 150020 65486
rect 150084 61130 150112 75140
rect 150176 72865 150204 75140
rect 150162 72856 150218 72865
rect 150162 72791 150218 72800
rect 150268 72282 150296 75140
rect 150360 72729 150388 75140
rect 150452 73234 150480 75140
rect 150440 73228 150492 73234
rect 150440 73170 150492 73176
rect 150438 73128 150494 73137
rect 150438 73063 150494 73072
rect 150346 72720 150402 72729
rect 150346 72655 150402 72664
rect 150452 72622 150480 73063
rect 150440 72616 150492 72622
rect 150440 72558 150492 72564
rect 150256 72276 150308 72282
rect 150256 72218 150308 72224
rect 150544 65686 150572 75140
rect 150164 65680 150216 65686
rect 150164 65622 150216 65628
rect 150532 65680 150584 65686
rect 150532 65622 150584 65628
rect 150072 61124 150124 61130
rect 150072 61066 150124 61072
rect 150176 60734 150204 65622
rect 150532 65544 150584 65550
rect 150532 65486 150584 65492
rect 150084 60706 150204 60734
rect 149980 42220 150032 42226
rect 149980 42162 150032 42168
rect 150084 31278 150112 60706
rect 150072 31272 150124 31278
rect 150072 31214 150124 31220
rect 149704 27124 149756 27130
rect 149704 27066 149756 27072
rect 150544 15978 150572 65486
rect 150636 61470 150664 75140
rect 150624 61464 150676 61470
rect 150624 61406 150676 61412
rect 150728 16046 150756 75140
rect 150820 67590 150848 75140
rect 150808 67584 150860 67590
rect 150808 67526 150860 67532
rect 150912 65362 150940 75140
rect 151004 65550 151032 75140
rect 151096 72758 151124 75140
rect 151084 72752 151136 72758
rect 151084 72694 151136 72700
rect 151082 72448 151138 72457
rect 151082 72383 151138 72392
rect 151096 71913 151124 72383
rect 151082 71904 151138 71913
rect 151082 71839 151138 71848
rect 150992 65544 151044 65550
rect 150992 65486 151044 65492
rect 151188 65482 151216 75140
rect 151280 70106 151308 75140
rect 151372 73234 151400 75140
rect 151360 73228 151412 73234
rect 151360 73170 151412 73176
rect 151360 72752 151412 72758
rect 151360 72694 151412 72700
rect 151268 70100 151320 70106
rect 151268 70042 151320 70048
rect 151268 65680 151320 65686
rect 151268 65622 151320 65628
rect 151176 65476 151228 65482
rect 151176 65418 151228 65424
rect 150912 65334 151216 65362
rect 151084 65272 151136 65278
rect 151084 65214 151136 65220
rect 151096 60042 151124 65214
rect 151084 60036 151136 60042
rect 151084 59978 151136 59984
rect 151188 51882 151216 65334
rect 151176 51876 151228 51882
rect 151176 51818 151228 51824
rect 151280 28490 151308 65622
rect 151268 28484 151320 28490
rect 151268 28426 151320 28432
rect 151372 27062 151400 72694
rect 151464 72593 151492 75140
rect 151556 72729 151584 75140
rect 151648 73953 151676 75140
rect 151634 73944 151690 73953
rect 151634 73879 151690 73888
rect 151636 72752 151688 72758
rect 151542 72720 151598 72729
rect 151636 72694 151688 72700
rect 151542 72655 151598 72664
rect 151450 72584 151506 72593
rect 151450 72519 151506 72528
rect 151648 70394 151676 72694
rect 151740 72457 151768 75140
rect 151726 72448 151782 72457
rect 151726 72383 151782 72392
rect 151464 70366 151676 70394
rect 151360 27056 151412 27062
rect 151360 26998 151412 27004
rect 151464 25702 151492 70366
rect 151544 67584 151596 67590
rect 151544 67526 151596 67532
rect 151452 25696 151504 25702
rect 151452 25638 151504 25644
rect 151556 18698 151584 67526
rect 151832 65550 151860 75140
rect 151924 71942 151952 75140
rect 151912 71936 151964 71942
rect 151912 71878 151964 71884
rect 152016 71330 152044 75140
rect 152004 71324 152056 71330
rect 152004 71266 152056 71272
rect 151820 65544 151872 65550
rect 151820 65486 151872 65492
rect 152108 60734 152136 75140
rect 152200 72418 152228 75140
rect 152292 74633 152320 75140
rect 152278 74624 152334 74633
rect 152278 74559 152334 74568
rect 152280 74180 152332 74186
rect 152280 74122 152332 74128
rect 152292 73302 152320 74122
rect 152280 73296 152332 73302
rect 152280 73238 152332 73244
rect 152280 73160 152332 73166
rect 152280 73102 152332 73108
rect 152188 72412 152240 72418
rect 152188 72354 152240 72360
rect 152188 72276 152240 72282
rect 152188 72218 152240 72224
rect 152200 66910 152228 72218
rect 152188 66904 152240 66910
rect 152188 66846 152240 66852
rect 152292 64138 152320 73102
rect 152384 73030 152412 75140
rect 152372 73024 152424 73030
rect 152372 72966 152424 72972
rect 152372 72820 152424 72826
rect 152372 72762 152424 72768
rect 152384 64258 152412 72762
rect 152476 64258 152504 75140
rect 152568 72706 152596 75140
rect 152660 72826 152688 75140
rect 152752 74186 152780 75140
rect 152740 74180 152792 74186
rect 152740 74122 152792 74128
rect 152740 73976 152792 73982
rect 152740 73918 152792 73924
rect 152752 72865 152780 73918
rect 152738 72856 152794 72865
rect 152648 72820 152700 72826
rect 152738 72791 152794 72800
rect 152648 72762 152700 72768
rect 152568 72678 152780 72706
rect 152648 72616 152700 72622
rect 152648 72558 152700 72564
rect 152660 69222 152688 72558
rect 152648 69216 152700 69222
rect 152648 69158 152700 69164
rect 152372 64252 152424 64258
rect 152372 64194 152424 64200
rect 152464 64252 152516 64258
rect 152464 64194 152516 64200
rect 152292 64110 152504 64138
rect 152372 64048 152424 64054
rect 152372 63990 152424 63996
rect 152108 60706 152228 60734
rect 151544 18692 151596 18698
rect 151544 18634 151596 18640
rect 151084 17264 151136 17270
rect 151084 17206 151136 17212
rect 150716 16040 150768 16046
rect 150716 15982 150768 15988
rect 150532 15972 150584 15978
rect 150532 15914 150584 15920
rect 149428 9172 149480 9178
rect 149428 9114 149480 9120
rect 151096 4010 151124 17206
rect 152200 15910 152228 60706
rect 152188 15904 152240 15910
rect 151174 15872 151230 15881
rect 152188 15846 152240 15852
rect 151174 15807 151230 15816
rect 151084 4004 151136 4010
rect 151084 3946 151136 3952
rect 151188 3670 151216 15807
rect 151820 6180 151872 6186
rect 151820 6122 151872 6128
rect 149520 3664 149572 3670
rect 149520 3606 149572 3612
rect 151176 3664 151228 3670
rect 151176 3606 151228 3612
rect 149532 480 149560 3606
rect 150624 3596 150676 3602
rect 150624 3538 150676 3544
rect 150636 480 150664 3538
rect 151832 480 151860 6122
rect 152384 4894 152412 63990
rect 152476 58886 152504 64110
rect 152464 58880 152516 58886
rect 152464 58822 152516 58828
rect 152752 45014 152780 72678
rect 152740 45008 152792 45014
rect 152740 44950 152792 44956
rect 152844 42158 152872 75140
rect 152936 72622 152964 75140
rect 153028 72729 153056 75140
rect 153120 73982 153148 75140
rect 153108 73976 153160 73982
rect 153108 73918 153160 73924
rect 153106 73536 153162 73545
rect 153106 73471 153162 73480
rect 153120 73001 153148 73471
rect 153106 72992 153162 73001
rect 153106 72927 153162 72936
rect 153108 72888 153160 72894
rect 153108 72830 153160 72836
rect 153014 72720 153070 72729
rect 153014 72655 153070 72664
rect 153120 72622 153148 72830
rect 152924 72616 152976 72622
rect 152924 72558 152976 72564
rect 153108 72616 153160 72622
rect 153108 72558 153160 72564
rect 153212 69970 153240 75140
rect 153304 73166 153332 75140
rect 153292 73160 153344 73166
rect 153292 73102 153344 73108
rect 153290 72992 153346 73001
rect 153290 72927 153346 72936
rect 153304 72486 153332 72927
rect 153292 72480 153344 72486
rect 153292 72422 153344 72428
rect 153292 72344 153344 72350
rect 153292 72286 153344 72292
rect 153200 69964 153252 69970
rect 153200 69906 153252 69912
rect 153200 65612 153252 65618
rect 153200 65554 153252 65560
rect 152924 65544 152976 65550
rect 152924 65486 152976 65492
rect 152832 42152 152884 42158
rect 152832 42094 152884 42100
rect 152936 24342 152964 65486
rect 152924 24336 152976 24342
rect 152924 24278 152976 24284
rect 153212 6390 153240 65554
rect 153304 60734 153332 72286
rect 153396 65226 153424 75140
rect 153488 65482 153516 75140
rect 153580 65686 153608 75140
rect 153568 65680 153620 65686
rect 153568 65622 153620 65628
rect 153476 65476 153528 65482
rect 153476 65418 153528 65424
rect 153672 65362 153700 75140
rect 153764 65550 153792 75140
rect 153856 72826 153884 75140
rect 153844 72820 153896 72826
rect 153844 72762 153896 72768
rect 153844 72548 153896 72554
rect 153844 72490 153896 72496
rect 153856 72321 153884 72490
rect 153842 72312 153898 72321
rect 153842 72247 153898 72256
rect 153752 65544 153804 65550
rect 153752 65486 153804 65492
rect 153948 65498 153976 75140
rect 154040 65618 154068 75140
rect 154132 72457 154160 75140
rect 154224 72865 154252 75140
rect 154210 72856 154266 72865
rect 154210 72791 154266 72800
rect 154316 72729 154344 75140
rect 154302 72720 154358 72729
rect 154302 72655 154358 72664
rect 154118 72448 154174 72457
rect 154118 72383 154174 72392
rect 154408 72010 154436 75140
rect 154500 72593 154528 75140
rect 154486 72584 154542 72593
rect 154486 72519 154542 72528
rect 154488 72208 154540 72214
rect 154488 72150 154540 72156
rect 154396 72004 154448 72010
rect 154396 71946 154448 71952
rect 154500 66978 154528 72150
rect 154488 66972 154540 66978
rect 154488 66914 154540 66920
rect 154396 65680 154448 65686
rect 154396 65622 154448 65628
rect 154028 65612 154080 65618
rect 154028 65554 154080 65560
rect 154212 65544 154264 65550
rect 153948 65470 154160 65498
rect 154212 65486 154264 65492
rect 153672 65334 154068 65362
rect 153396 65198 153976 65226
rect 153304 60706 153884 60734
rect 153856 38010 153884 60706
rect 153948 58818 153976 65198
rect 153936 58812 153988 58818
rect 153936 58754 153988 58760
rect 154040 53310 154068 65334
rect 154028 53304 154080 53310
rect 154028 53246 154080 53252
rect 154132 47666 154160 65470
rect 154120 47660 154172 47666
rect 154120 47602 154172 47608
rect 153844 38004 153896 38010
rect 153844 37946 153896 37952
rect 154224 14482 154252 65486
rect 154304 65476 154356 65482
rect 154304 65418 154356 65424
rect 154212 14476 154264 14482
rect 154212 14418 154264 14424
rect 154316 13258 154344 65418
rect 154304 13252 154356 13258
rect 154304 13194 154356 13200
rect 153844 13116 153896 13122
rect 153844 13058 153896 13064
rect 153200 6384 153252 6390
rect 153200 6326 153252 6332
rect 152372 4888 152424 4894
rect 152372 4830 152424 4836
rect 153016 4004 153068 4010
rect 153016 3946 153068 3952
rect 153028 480 153056 3946
rect 153856 3330 153884 13058
rect 154408 9110 154436 65622
rect 154592 65278 154620 75140
rect 154684 72622 154712 75140
rect 154672 72616 154724 72622
rect 154672 72558 154724 72564
rect 154672 65612 154724 65618
rect 154672 65554 154724 65560
rect 154580 65272 154632 65278
rect 154580 65214 154632 65220
rect 154396 9104 154448 9110
rect 154396 9046 154448 9052
rect 154684 6322 154712 65554
rect 154776 60734 154804 75140
rect 154868 72706 154896 75140
rect 154960 73166 154988 75140
rect 154948 73160 155000 73166
rect 154948 73102 155000 73108
rect 154868 72678 154988 72706
rect 154856 72616 154908 72622
rect 154856 72558 154908 72564
rect 154868 65346 154896 72558
rect 154960 65890 154988 72678
rect 154948 65884 155000 65890
rect 154948 65826 155000 65832
rect 155052 65498 155080 75140
rect 155144 65686 155172 75140
rect 155132 65680 155184 65686
rect 155132 65622 155184 65628
rect 155236 65618 155264 75140
rect 155224 65612 155276 65618
rect 155224 65554 155276 65560
rect 155052 65470 155264 65498
rect 154856 65340 154908 65346
rect 154856 65282 154908 65288
rect 154776 60706 155172 60734
rect 155144 54602 155172 60706
rect 155132 54596 155184 54602
rect 155132 54538 155184 54544
rect 155236 50454 155264 65470
rect 155224 50448 155276 50454
rect 155224 50390 155276 50396
rect 155328 43586 155356 75140
rect 155420 65498 155448 75140
rect 155512 73098 155540 75140
rect 155500 73092 155552 73098
rect 155500 73034 155552 73040
rect 155604 72865 155632 75140
rect 155590 72856 155646 72865
rect 155500 72820 155552 72826
rect 155590 72791 155646 72800
rect 155500 72762 155552 72768
rect 155512 72214 155540 72762
rect 155696 72593 155724 75140
rect 155788 72729 155816 75140
rect 155774 72720 155830 72729
rect 155774 72655 155830 72664
rect 155682 72584 155738 72593
rect 155682 72519 155738 72528
rect 155880 72457 155908 75140
rect 155866 72448 155922 72457
rect 155866 72383 155922 72392
rect 155500 72208 155552 72214
rect 155500 72150 155552 72156
rect 155500 71732 155552 71738
rect 155500 71674 155552 71680
rect 155512 70174 155540 71674
rect 155500 70168 155552 70174
rect 155500 70110 155552 70116
rect 155972 67522 156000 75140
rect 156064 73098 156092 75140
rect 156052 73092 156104 73098
rect 156052 73034 156104 73040
rect 156156 72622 156184 75140
rect 156144 72616 156196 72622
rect 156144 72558 156196 72564
rect 156142 72312 156198 72321
rect 156142 72247 156144 72256
rect 156196 72247 156198 72256
rect 156144 72218 156196 72224
rect 155960 67516 156012 67522
rect 155960 67458 156012 67464
rect 155776 65884 155828 65890
rect 155776 65826 155828 65832
rect 155420 65470 155724 65498
rect 155408 65408 155460 65414
rect 155408 65350 155460 65356
rect 155316 43580 155368 43586
rect 155316 43522 155368 43528
rect 155222 38040 155278 38049
rect 155222 37975 155278 37984
rect 154672 6316 154724 6322
rect 154672 6258 154724 6264
rect 155236 3534 155264 37975
rect 155420 36582 155448 65350
rect 155592 65340 155644 65346
rect 155592 65282 155644 65288
rect 155500 65272 155552 65278
rect 155500 65214 155552 65220
rect 155408 36576 155460 36582
rect 155408 36518 155460 36524
rect 155512 33862 155540 65214
rect 155500 33856 155552 33862
rect 155500 33798 155552 33804
rect 155604 13190 155632 65282
rect 155592 13184 155644 13190
rect 155592 13126 155644 13132
rect 155696 10470 155724 65470
rect 155684 10464 155736 10470
rect 155684 10406 155736 10412
rect 155788 7682 155816 65826
rect 156248 65686 156276 75140
rect 156340 71806 156368 75140
rect 156328 71800 156380 71806
rect 156328 71742 156380 71748
rect 156432 71194 156460 75140
rect 156420 71188 156472 71194
rect 156420 71130 156472 71136
rect 156524 70394 156552 75140
rect 156616 72350 156644 75140
rect 156604 72344 156656 72350
rect 156604 72286 156656 72292
rect 156708 70394 156736 75140
rect 156340 70366 156552 70394
rect 156616 70366 156736 70394
rect 156236 65680 156288 65686
rect 156236 65622 156288 65628
rect 156340 64002 156368 70366
rect 155972 63974 156368 64002
rect 155972 28422 156000 63974
rect 156616 63458 156644 70366
rect 156800 67674 156828 75140
rect 156892 71890 156920 75140
rect 156984 72026 157012 75140
rect 157076 72162 157104 75140
rect 157168 72962 157196 75140
rect 157156 72956 157208 72962
rect 157156 72898 157208 72904
rect 157260 72593 157288 75140
rect 157246 72584 157302 72593
rect 157246 72519 157302 72528
rect 157248 72480 157300 72486
rect 157248 72422 157300 72428
rect 157076 72134 157196 72162
rect 156984 71998 157104 72026
rect 156892 71862 157012 71890
rect 156880 71800 156932 71806
rect 156880 71742 156932 71748
rect 156248 63430 156644 63458
rect 156708 67646 156828 67674
rect 155960 28416 156012 28422
rect 155960 28358 156012 28364
rect 155776 7676 155828 7682
rect 155776 7618 155828 7624
rect 156248 3806 156276 63430
rect 156420 63368 156472 63374
rect 156420 63310 156472 63316
rect 156236 3800 156288 3806
rect 156236 3742 156288 3748
rect 156432 3670 156460 63310
rect 156708 61402 156736 67646
rect 156788 67516 156840 67522
rect 156788 67458 156840 67464
rect 156696 61396 156748 61402
rect 156696 61338 156748 61344
rect 156800 47598 156828 67458
rect 156788 47592 156840 47598
rect 156788 47534 156840 47540
rect 156892 44946 156920 71742
rect 156880 44940 156932 44946
rect 156880 44882 156932 44888
rect 156602 42120 156658 42129
rect 156602 42055 156658 42064
rect 155408 3664 155460 3670
rect 155408 3606 155460 3612
rect 156420 3664 156472 3670
rect 156420 3606 156472 3612
rect 154212 3528 154264 3534
rect 154212 3470 154264 3476
rect 155224 3528 155276 3534
rect 155224 3470 155276 3476
rect 153844 3324 153896 3330
rect 153844 3266 153896 3272
rect 154224 480 154252 3470
rect 155420 480 155448 3606
rect 156616 480 156644 42055
rect 156696 36644 156748 36650
rect 156696 36586 156748 36592
rect 156708 3602 156736 36586
rect 156984 29714 157012 71862
rect 157076 63374 157104 71998
rect 157168 71913 157196 72134
rect 157154 71904 157210 71913
rect 157154 71839 157210 71848
rect 157260 70038 157288 72422
rect 157248 70032 157300 70038
rect 157248 69974 157300 69980
rect 157064 63368 157116 63374
rect 157064 63310 157116 63316
rect 156972 29708 157024 29714
rect 156972 29650 157024 29656
rect 157352 29646 157380 75140
rect 157444 68610 157472 75140
rect 157536 73137 157564 75140
rect 157522 73128 157578 73137
rect 157522 73063 157578 73072
rect 157524 72820 157576 72826
rect 157524 72762 157576 72768
rect 157536 71874 157564 72762
rect 157524 71868 157576 71874
rect 157524 71810 157576 71816
rect 157432 68604 157484 68610
rect 157432 68546 157484 68552
rect 157432 65544 157484 65550
rect 157432 65486 157484 65492
rect 157340 29640 157392 29646
rect 157340 29582 157392 29588
rect 157444 17338 157472 65486
rect 157628 17406 157656 75140
rect 157720 74905 157748 75140
rect 157706 74896 157762 74905
rect 157706 74831 157762 74840
rect 157708 74792 157760 74798
rect 157708 74734 157760 74740
rect 157720 73273 157748 74734
rect 157706 73264 157762 73273
rect 157706 73199 157762 73208
rect 157708 73160 157760 73166
rect 157708 73102 157760 73108
rect 157720 72418 157748 73102
rect 157708 72412 157760 72418
rect 157708 72354 157760 72360
rect 157708 71800 157760 71806
rect 157708 71742 157760 71748
rect 157720 61198 157748 71742
rect 157812 69834 157840 75140
rect 157800 69828 157852 69834
rect 157800 69770 157852 69776
rect 157904 65550 157932 75140
rect 157996 73234 158024 75140
rect 157984 73228 158036 73234
rect 157984 73170 158036 73176
rect 157982 73128 158038 73137
rect 157982 73063 158038 73072
rect 157996 72729 158024 73063
rect 157982 72720 158038 72729
rect 157982 72655 158038 72664
rect 157982 72176 158038 72185
rect 157982 72111 158038 72120
rect 157996 70718 158024 72111
rect 157984 70712 158036 70718
rect 157984 70654 158036 70660
rect 158088 69766 158116 75140
rect 158076 69760 158128 69766
rect 158076 69702 158128 69708
rect 157892 65544 157944 65550
rect 157892 65486 157944 65492
rect 158180 61282 158208 75140
rect 158272 72298 158300 75140
rect 158364 72729 158392 75140
rect 158350 72720 158406 72729
rect 158350 72655 158406 72664
rect 158456 72457 158484 75140
rect 158548 72729 158576 75140
rect 158534 72720 158590 72729
rect 158534 72655 158590 72664
rect 158640 72593 158668 75140
rect 158626 72584 158682 72593
rect 158626 72519 158682 72528
rect 158442 72448 158498 72457
rect 158442 72383 158498 72392
rect 158626 72448 158682 72457
rect 158626 72383 158682 72392
rect 158272 72270 158392 72298
rect 158640 72282 158668 72383
rect 158364 72185 158392 72270
rect 158628 72276 158680 72282
rect 158628 72218 158680 72224
rect 158350 72176 158406 72185
rect 158260 72140 158312 72146
rect 158350 72111 158406 72120
rect 158260 72082 158312 72088
rect 158272 62898 158300 72082
rect 158732 65550 158760 75140
rect 158824 73302 158852 75140
rect 158916 73817 158944 75140
rect 158902 73808 158958 73817
rect 158902 73743 158958 73752
rect 158902 73400 158958 73409
rect 158902 73335 158904 73344
rect 158956 73335 158958 73344
rect 158904 73306 158956 73312
rect 158812 73296 158864 73302
rect 158812 73238 158864 73244
rect 158812 73160 158864 73166
rect 158812 73102 158864 73108
rect 158720 65544 158772 65550
rect 158720 65486 158772 65492
rect 158824 65142 158852 73102
rect 158904 73092 158956 73098
rect 158904 73034 158956 73040
rect 158916 71942 158944 73034
rect 158904 71936 158956 71942
rect 158904 71878 158956 71884
rect 158904 71800 158956 71806
rect 158904 71742 158956 71748
rect 158916 65278 158944 71742
rect 158904 65272 158956 65278
rect 158904 65214 158956 65220
rect 159008 65210 159036 75140
rect 158996 65204 159048 65210
rect 158996 65146 159048 65152
rect 158812 65136 158864 65142
rect 158812 65078 158864 65084
rect 158260 62892 158312 62898
rect 158260 62834 158312 62840
rect 157812 61254 158208 61282
rect 157708 61192 157760 61198
rect 157708 61134 157760 61140
rect 157616 17400 157668 17406
rect 157616 17342 157668 17348
rect 157432 17332 157484 17338
rect 157432 17274 157484 17280
rect 157812 17270 157840 61254
rect 157984 61192 158036 61198
rect 157984 61134 158036 61140
rect 157800 17264 157852 17270
rect 157800 17206 157852 17212
rect 157996 4962 158024 61134
rect 159100 60734 159128 75140
rect 159192 74186 159220 75140
rect 159180 74180 159232 74186
rect 159180 74122 159232 74128
rect 159180 73092 159232 73098
rect 159180 73034 159232 73040
rect 159192 72729 159220 73034
rect 159178 72720 159234 72729
rect 159178 72655 159234 72664
rect 159180 65544 159232 65550
rect 159180 65486 159232 65492
rect 159008 60706 159128 60734
rect 158076 29776 158128 29782
rect 158076 29718 158128 29724
rect 157984 4956 158036 4962
rect 157984 4898 158036 4904
rect 156696 3596 156748 3602
rect 156696 3538 156748 3544
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 157812 480 157840 3470
rect 158088 2990 158116 29718
rect 159008 11762 159036 60706
rect 158996 11756 159048 11762
rect 158996 11698 159048 11704
rect 159192 9042 159220 65486
rect 159284 65414 159312 75140
rect 159272 65408 159324 65414
rect 159272 65350 159324 65356
rect 159376 65362 159404 75140
rect 159468 72826 159496 75140
rect 159456 72820 159508 72826
rect 159456 72762 159508 72768
rect 159560 65498 159588 75140
rect 159652 72729 159680 75140
rect 159638 72720 159694 72729
rect 159638 72655 159694 72664
rect 159744 65890 159772 75140
rect 159836 72593 159864 75140
rect 159928 72729 159956 75140
rect 160020 73098 160048 75140
rect 160008 73092 160060 73098
rect 160008 73034 160060 73040
rect 160008 72820 160060 72826
rect 160008 72762 160060 72768
rect 159914 72720 159970 72729
rect 159914 72655 159970 72664
rect 159822 72584 159878 72593
rect 159822 72519 159878 72528
rect 159732 65884 159784 65890
rect 159732 65826 159784 65832
rect 159560 65470 159864 65498
rect 160020 65482 160048 72762
rect 160112 65618 160140 75140
rect 160204 69698 160232 75140
rect 160296 72826 160324 75140
rect 160284 72820 160336 72826
rect 160284 72762 160336 72768
rect 160282 72720 160338 72729
rect 160282 72655 160338 72664
rect 160296 70394 160324 72655
rect 160388 72078 160416 75140
rect 160376 72072 160428 72078
rect 160376 72014 160428 72020
rect 160296 70366 160416 70394
rect 160192 69692 160244 69698
rect 160192 69634 160244 69640
rect 160100 65612 160152 65618
rect 160100 65554 160152 65560
rect 159732 65408 159784 65414
rect 159376 65334 159680 65362
rect 159732 65350 159784 65356
rect 159364 65272 159416 65278
rect 159364 65214 159416 65220
rect 159376 20058 159404 65214
rect 159548 65204 159600 65210
rect 159548 65146 159600 65152
rect 159456 65136 159508 65142
rect 159456 65078 159508 65084
rect 159468 54534 159496 65078
rect 159456 54528 159508 54534
rect 159456 54470 159508 54476
rect 159560 43518 159588 65146
rect 159548 43512 159600 43518
rect 159548 43454 159600 43460
rect 159652 40798 159680 65334
rect 159640 40792 159692 40798
rect 159640 40734 159692 40740
rect 159744 31210 159772 65350
rect 159732 31204 159784 31210
rect 159732 31146 159784 31152
rect 159836 28354 159864 65470
rect 160008 65476 160060 65482
rect 160008 65418 160060 65424
rect 159824 28348 159876 28354
rect 159824 28290 159876 28296
rect 160388 26994 160416 70366
rect 160480 65550 160508 75140
rect 160572 72457 160600 75140
rect 160558 72448 160614 72457
rect 160558 72383 160614 72392
rect 160664 70394 160692 75140
rect 160756 72944 160784 75140
rect 160848 73234 160876 75140
rect 160836 73228 160888 73234
rect 160836 73170 160888 73176
rect 160756 72916 160876 72944
rect 160744 72820 160796 72826
rect 160744 72762 160796 72768
rect 160756 71806 160784 72762
rect 160848 72486 160876 72916
rect 160836 72480 160888 72486
rect 160836 72422 160888 72428
rect 160940 72282 160968 75140
rect 161032 72729 161060 75140
rect 161124 72944 161152 75140
rect 161216 73545 161244 75140
rect 161202 73536 161258 73545
rect 161202 73471 161258 73480
rect 161308 73273 161336 75140
rect 161294 73264 161350 73273
rect 161294 73199 161350 73208
rect 161124 72916 161336 72944
rect 161018 72720 161074 72729
rect 161018 72655 161074 72664
rect 160928 72276 160980 72282
rect 160928 72218 160980 72224
rect 161204 72276 161256 72282
rect 161204 72218 161256 72224
rect 160928 72072 160980 72078
rect 160928 72014 160980 72020
rect 160744 71800 160796 71806
rect 160744 71742 160796 71748
rect 160742 71360 160798 71369
rect 160742 71295 160798 71304
rect 160572 70366 160692 70394
rect 160468 65544 160520 65550
rect 160468 65486 160520 65492
rect 160572 60734 160600 70366
rect 160756 60734 160784 71295
rect 160836 65544 160888 65550
rect 160836 65486 160888 65492
rect 160480 60706 160600 60734
rect 160664 60706 160784 60734
rect 160376 26988 160428 26994
rect 160376 26930 160428 26936
rect 160480 25634 160508 60706
rect 160468 25628 160520 25634
rect 160468 25570 160520 25576
rect 160664 24206 160692 60706
rect 160848 44878 160876 65486
rect 160836 44872 160888 44878
rect 160836 44814 160888 44820
rect 160940 40730 160968 72014
rect 161216 67634 161244 72218
rect 161032 67606 161244 67634
rect 160744 40724 160796 40730
rect 160744 40666 160796 40672
rect 160928 40724 160980 40730
rect 160928 40666 160980 40672
rect 160652 24200 160704 24206
rect 160652 24142 160704 24148
rect 159364 20052 159416 20058
rect 159364 19994 159416 20000
rect 159180 9036 159232 9042
rect 159180 8978 159232 8984
rect 160756 4010 160784 40666
rect 161032 39438 161060 67606
rect 161308 67182 161336 72916
rect 161400 72593 161428 75140
rect 161386 72584 161442 72593
rect 161386 72519 161442 72528
rect 161388 72480 161440 72486
rect 161388 72422 161440 72428
rect 161400 71194 161428 72422
rect 161388 71188 161440 71194
rect 161388 71130 161440 71136
rect 161296 67176 161348 67182
rect 161296 67118 161348 67124
rect 161112 65612 161164 65618
rect 161112 65554 161164 65560
rect 161020 39432 161072 39438
rect 161020 39374 161072 39380
rect 161124 35222 161152 65554
rect 161112 35216 161164 35222
rect 161112 35158 161164 35164
rect 161492 22778 161520 75140
rect 161584 72706 161612 75140
rect 161676 73778 161704 75140
rect 161664 73772 161716 73778
rect 161664 73714 161716 73720
rect 161584 72678 161704 72706
rect 161676 65278 161704 72678
rect 161768 70394 161796 75140
rect 161860 72554 161888 75140
rect 161848 72548 161900 72554
rect 161848 72490 161900 72496
rect 161952 72486 161980 75140
rect 161940 72480 161992 72486
rect 161940 72422 161992 72428
rect 161940 72208 161992 72214
rect 161940 72150 161992 72156
rect 161952 71874 161980 72150
rect 161940 71868 161992 71874
rect 161940 71810 161992 71816
rect 161768 70366 161888 70394
rect 161664 65272 161716 65278
rect 161664 65214 161716 65220
rect 161860 63510 161888 70366
rect 161940 69964 161992 69970
rect 161940 69906 161992 69912
rect 161952 69222 161980 69906
rect 161940 69216 161992 69222
rect 161940 69158 161992 69164
rect 162044 65618 162072 75140
rect 162032 65612 162084 65618
rect 162032 65554 162084 65560
rect 162136 65498 162164 75140
rect 162228 70417 162256 75140
rect 162214 70408 162270 70417
rect 162214 70343 162270 70352
rect 162216 70304 162268 70310
rect 162216 70246 162268 70252
rect 162228 69290 162256 70246
rect 162216 69284 162268 69290
rect 162216 69226 162268 69232
rect 161952 65470 162164 65498
rect 161848 63504 161900 63510
rect 161848 63446 161900 63452
rect 161952 60734 161980 65470
rect 162320 65362 162348 75140
rect 161768 60706 161980 60734
rect 162136 65334 162348 65362
rect 161768 25566 161796 60706
rect 162136 51746 162164 65334
rect 162216 65272 162268 65278
rect 162216 65214 162268 65220
rect 162124 51740 162176 51746
rect 162124 51682 162176 51688
rect 162228 43450 162256 65214
rect 162412 63594 162440 75140
rect 162504 72593 162532 75140
rect 162596 73137 162624 75140
rect 162582 73128 162638 73137
rect 162582 73063 162638 73072
rect 162584 72888 162636 72894
rect 162584 72830 162636 72836
rect 162596 72758 162624 72830
rect 162584 72752 162636 72758
rect 162688 72729 162716 75140
rect 162584 72694 162636 72700
rect 162674 72720 162730 72729
rect 162674 72655 162730 72664
rect 162490 72584 162546 72593
rect 162490 72519 162546 72528
rect 162584 72548 162636 72554
rect 162584 72490 162636 72496
rect 162492 65612 162544 65618
rect 162492 65554 162544 65560
rect 162320 63566 162440 63594
rect 162216 43444 162268 43450
rect 162216 43386 162268 43392
rect 162320 42090 162348 63566
rect 162400 63504 162452 63510
rect 162400 63446 162452 63452
rect 162308 42084 162360 42090
rect 162308 42026 162360 42032
rect 162412 33794 162440 63446
rect 162400 33788 162452 33794
rect 162400 33730 162452 33736
rect 162504 32434 162532 65554
rect 162596 32502 162624 72490
rect 162676 72480 162728 72486
rect 162780 72457 162808 75140
rect 162676 72422 162728 72428
rect 162766 72448 162822 72457
rect 162688 64190 162716 72422
rect 162766 72383 162822 72392
rect 162766 70408 162822 70417
rect 162766 70343 162822 70352
rect 162676 64184 162728 64190
rect 162676 64126 162728 64132
rect 162780 62830 162808 70343
rect 162872 65550 162900 75140
rect 162860 65544 162912 65550
rect 162860 65486 162912 65492
rect 162964 65278 162992 75140
rect 163056 74050 163084 75140
rect 163044 74044 163096 74050
rect 163044 73986 163096 73992
rect 163044 73364 163096 73370
rect 163044 73306 163096 73312
rect 163056 72214 163084 73306
rect 163148 72486 163176 75140
rect 163136 72480 163188 72486
rect 163136 72422 163188 72428
rect 163044 72208 163096 72214
rect 163044 72150 163096 72156
rect 163240 70394 163268 75140
rect 163332 73914 163360 75140
rect 163320 73908 163372 73914
rect 163320 73850 163372 73856
rect 163424 72842 163452 75140
rect 163332 72814 163452 72842
rect 163332 71913 163360 72814
rect 163412 72548 163464 72554
rect 163412 72490 163464 72496
rect 163318 71904 163374 71913
rect 163318 71839 163374 71848
rect 163240 70366 163360 70394
rect 163228 65612 163280 65618
rect 163228 65554 163280 65560
rect 162952 65272 163004 65278
rect 162952 65214 163004 65220
rect 162768 62824 162820 62830
rect 162768 62766 162820 62772
rect 162584 32496 162636 32502
rect 162584 32438 162636 32444
rect 162492 32428 162544 32434
rect 162492 32370 162544 32376
rect 162124 31068 162176 31074
rect 162124 31010 162176 31016
rect 161756 25560 161808 25566
rect 161756 25502 161808 25508
rect 161480 22772 161532 22778
rect 161480 22714 161532 22720
rect 160744 4004 160796 4010
rect 160744 3946 160796 3952
rect 161294 3904 161350 3913
rect 161294 3839 161350 3848
rect 158904 3324 158956 3330
rect 158904 3266 158956 3272
rect 158076 2984 158128 2990
rect 158076 2926 158128 2932
rect 158916 480 158944 3266
rect 160100 2984 160152 2990
rect 160100 2926 160152 2932
rect 160112 480 160140 2926
rect 161308 480 161336 3839
rect 162136 3534 162164 31010
rect 163240 7614 163268 65554
rect 163332 65346 163360 70366
rect 163424 65498 163452 72490
rect 163516 70394 163544 75140
rect 163608 72554 163636 75140
rect 163596 72548 163648 72554
rect 163596 72490 163648 72496
rect 163516 70366 163636 70394
rect 163424 65470 163544 65498
rect 163412 65408 163464 65414
rect 163412 65350 163464 65356
rect 163320 65340 163372 65346
rect 163320 65282 163372 65288
rect 163424 58750 163452 65350
rect 163412 58744 163464 58750
rect 163412 58686 163464 58692
rect 163516 57254 163544 65470
rect 163504 57248 163556 57254
rect 163504 57190 163556 57196
rect 163608 53242 163636 70366
rect 163700 65618 163728 75140
rect 163688 65612 163740 65618
rect 163688 65554 163740 65560
rect 163792 65498 163820 75140
rect 163700 65470 163820 65498
rect 163596 53236 163648 53242
rect 163596 53178 163648 53184
rect 163700 39370 163728 65470
rect 163884 65414 163912 75140
rect 163976 72593 164004 75140
rect 163962 72584 164018 72593
rect 163962 72519 164018 72528
rect 163964 72480 164016 72486
rect 164068 72457 164096 75140
rect 164160 72729 164188 75140
rect 164146 72720 164202 72729
rect 164146 72655 164202 72664
rect 164146 72584 164202 72593
rect 164146 72519 164202 72528
rect 163964 72422 164016 72428
rect 164054 72448 164110 72457
rect 163872 65408 163924 65414
rect 163872 65350 163924 65356
rect 163780 65340 163832 65346
rect 163780 65282 163832 65288
rect 163688 39364 163740 39370
rect 163688 39306 163740 39312
rect 163792 31142 163820 65282
rect 163872 65272 163924 65278
rect 163872 65214 163924 65220
rect 163780 31136 163832 31142
rect 163780 31078 163832 31084
rect 163884 24138 163912 65214
rect 163872 24132 163924 24138
rect 163872 24074 163924 24080
rect 163976 10334 164004 72422
rect 164054 72383 164110 72392
rect 164160 71058 164188 72519
rect 164148 71052 164200 71058
rect 164148 70994 164200 71000
rect 164252 65618 164280 75140
rect 164240 65612 164292 65618
rect 164240 65554 164292 65560
rect 164056 65544 164108 65550
rect 164056 65486 164108 65492
rect 163964 10328 164016 10334
rect 163964 10270 164016 10276
rect 164068 8974 164096 65486
rect 164344 65482 164372 75140
rect 164436 73982 164464 75140
rect 164424 73976 164476 73982
rect 164424 73918 164476 73924
rect 164424 73160 164476 73166
rect 164424 73102 164476 73108
rect 164436 72554 164464 73102
rect 164424 72548 164476 72554
rect 164424 72490 164476 72496
rect 164528 65550 164556 75140
rect 164620 72162 164648 75140
rect 164712 73846 164740 75140
rect 164700 73840 164752 73846
rect 164700 73782 164752 73788
rect 164620 72134 164740 72162
rect 164608 72072 164660 72078
rect 164608 72014 164660 72020
rect 164620 68474 164648 72014
rect 164712 68542 164740 72134
rect 164700 68536 164752 68542
rect 164700 68478 164752 68484
rect 164608 68468 164660 68474
rect 164608 68410 164660 68416
rect 164516 65544 164568 65550
rect 164516 65486 164568 65492
rect 164332 65476 164384 65482
rect 164332 65418 164384 65424
rect 164804 64546 164832 75140
rect 164620 64518 164832 64546
rect 164056 8968 164108 8974
rect 164056 8910 164108 8916
rect 163228 7608 163280 7614
rect 163228 7550 163280 7556
rect 164620 6254 164648 64518
rect 164896 60734 164924 75140
rect 164804 60706 164924 60734
rect 164608 6248 164660 6254
rect 164608 6190 164660 6196
rect 164804 6186 164832 60706
rect 164988 55894 165016 75140
rect 165080 71097 165108 75140
rect 165172 72078 165200 75140
rect 165160 72072 165212 72078
rect 165160 72014 165212 72020
rect 165066 71088 165122 71097
rect 165066 71023 165122 71032
rect 165264 70394 165292 75140
rect 165356 72729 165384 75140
rect 165342 72720 165398 72729
rect 165342 72655 165398 72664
rect 165448 72593 165476 75140
rect 165434 72584 165490 72593
rect 165434 72519 165490 72528
rect 165540 72457 165568 75140
rect 165526 72448 165582 72457
rect 165526 72383 165582 72392
rect 165632 71890 165660 75140
rect 165724 73098 165752 75140
rect 165712 73092 165764 73098
rect 165712 73034 165764 73040
rect 165710 72584 165766 72593
rect 165710 72519 165766 72528
rect 165724 72185 165752 72519
rect 165710 72176 165766 72185
rect 165710 72111 165766 72120
rect 165448 71862 165660 71890
rect 165710 71904 165766 71913
rect 165448 71346 165476 71862
rect 165710 71839 165766 71848
rect 165620 71800 165672 71806
rect 165620 71742 165672 71748
rect 165632 71618 165660 71742
rect 165724 71738 165752 71839
rect 165712 71732 165764 71738
rect 165712 71674 165764 71680
rect 165632 71590 165752 71618
rect 165448 71318 165660 71346
rect 165172 70366 165292 70394
rect 165068 65544 165120 65550
rect 165068 65486 165120 65492
rect 164976 55888 165028 55894
rect 164976 55830 165028 55836
rect 165080 53174 165108 65486
rect 165068 53168 165120 53174
rect 165068 53110 165120 53116
rect 165172 50386 165200 70366
rect 165632 65618 165660 71318
rect 165252 65612 165304 65618
rect 165252 65554 165304 65560
rect 165620 65612 165672 65618
rect 165620 65554 165672 65560
rect 165160 50380 165212 50386
rect 165160 50322 165212 50328
rect 165264 31074 165292 65554
rect 165344 65476 165396 65482
rect 165344 65418 165396 65424
rect 165252 31068 165304 31074
rect 165252 31010 165304 31016
rect 165356 13122 165384 65418
rect 165724 65414 165752 71590
rect 165816 65550 165844 75140
rect 165804 65544 165856 65550
rect 165804 65486 165856 65492
rect 165712 65408 165764 65414
rect 165712 65350 165764 65356
rect 165908 26926 165936 75140
rect 166000 60734 166028 75140
rect 166092 65498 166120 75140
rect 166184 65634 166212 75140
rect 166276 68338 166304 75140
rect 166368 72185 166396 75140
rect 166460 72457 166488 75140
rect 166552 72593 166580 75140
rect 166538 72584 166594 72593
rect 166538 72519 166594 72528
rect 166446 72448 166502 72457
rect 166446 72383 166502 72392
rect 166644 72185 166672 75140
rect 166354 72176 166410 72185
rect 166354 72111 166410 72120
rect 166630 72176 166686 72185
rect 166630 72111 166686 72120
rect 166736 72049 166764 75140
rect 166828 73545 166856 75140
rect 166814 73536 166870 73545
rect 166814 73471 166870 73480
rect 166920 73250 166948 75140
rect 166828 73222 166948 73250
rect 166828 72486 166856 73222
rect 166908 73092 166960 73098
rect 166908 73034 166960 73040
rect 166816 72480 166868 72486
rect 166816 72422 166868 72428
rect 166722 72040 166778 72049
rect 166722 71975 166778 71984
rect 166920 68406 166948 73034
rect 167012 72078 167040 75140
rect 167000 72072 167052 72078
rect 167000 72014 167052 72020
rect 167104 70786 167132 75140
rect 167196 71369 167224 75140
rect 167288 71505 167316 75140
rect 167380 72146 167408 75140
rect 167472 74458 167500 75140
rect 167564 74633 167592 75140
rect 167550 74624 167606 74633
rect 167550 74559 167606 74568
rect 167460 74452 167512 74458
rect 167460 74394 167512 74400
rect 167656 73574 167684 75140
rect 167748 74526 167776 75140
rect 167736 74520 167788 74526
rect 167736 74462 167788 74468
rect 167644 73568 167696 73574
rect 167644 73510 167696 73516
rect 167840 73098 167868 75140
rect 167932 73642 167960 75140
rect 167920 73636 167972 73642
rect 167920 73578 167972 73584
rect 167828 73092 167880 73098
rect 167828 73034 167880 73040
rect 168024 73030 168052 75140
rect 168116 73506 168144 75140
rect 168104 73500 168156 73506
rect 168104 73442 168156 73448
rect 167552 73024 167604 73030
rect 167552 72966 167604 72972
rect 168012 73024 168064 73030
rect 168012 72966 168064 72972
rect 167368 72140 167420 72146
rect 167368 72082 167420 72088
rect 167274 71496 167330 71505
rect 167274 71431 167330 71440
rect 167182 71360 167238 71369
rect 167182 71295 167238 71304
rect 167092 70780 167144 70786
rect 167092 70722 167144 70728
rect 167184 68876 167236 68882
rect 167184 68818 167236 68824
rect 166908 68400 166960 68406
rect 166908 68342 166960 68348
rect 166264 68332 166316 68338
rect 166264 68274 166316 68280
rect 166908 65884 166960 65890
rect 166908 65826 166960 65832
rect 166184 65606 166672 65634
rect 166540 65544 166592 65550
rect 166092 65470 166396 65498
rect 166540 65486 166592 65492
rect 166264 65408 166316 65414
rect 166264 65350 166316 65356
rect 166000 60706 166120 60734
rect 165896 26920 165948 26926
rect 165896 26862 165948 26868
rect 166092 18630 166120 60706
rect 166080 18624 166132 18630
rect 166080 18566 166132 18572
rect 165344 13116 165396 13122
rect 165344 13058 165396 13064
rect 164792 6180 164844 6186
rect 164792 6122 164844 6128
rect 166276 4826 166304 65350
rect 166368 60734 166396 65470
rect 166368 60706 166488 60734
rect 166460 58682 166488 60706
rect 166448 58676 166500 58682
rect 166448 58618 166500 58624
rect 166552 53106 166580 65486
rect 166540 53100 166592 53106
rect 166540 53042 166592 53048
rect 166644 37942 166672 65606
rect 166724 65612 166776 65618
rect 166724 65554 166776 65560
rect 166632 37936 166684 37942
rect 166632 37878 166684 37884
rect 166736 28286 166764 65554
rect 166920 65550 166948 65826
rect 166908 65544 166960 65550
rect 166908 65486 166960 65492
rect 166724 28280 166776 28286
rect 166724 28222 166776 28228
rect 166264 4820 166316 4826
rect 166264 4762 166316 4768
rect 162492 4004 162544 4010
rect 162492 3946 162544 3952
rect 162124 3528 162176 3534
rect 162124 3470 162176 3476
rect 162504 480 162532 3946
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 163700 480 163728 3470
rect 164896 480 164924 3538
rect 166080 3460 166132 3466
rect 166080 3402 166132 3408
rect 166092 480 166120 3402
rect 167196 480 167224 68818
rect 167564 51814 167592 72966
rect 167736 72820 167788 72826
rect 167736 72762 167788 72768
rect 167644 72684 167696 72690
rect 167644 72626 167696 72632
rect 167552 51808 167604 51814
rect 167552 51750 167604 51756
rect 167656 4010 167684 72626
rect 167748 71126 167776 72762
rect 168104 72752 168156 72758
rect 168104 72694 168156 72700
rect 167920 72004 167972 72010
rect 167920 71946 167972 71952
rect 167828 71868 167880 71874
rect 167828 71810 167880 71816
rect 167736 71120 167788 71126
rect 167736 71062 167788 71068
rect 167736 70712 167788 70718
rect 167736 70654 167788 70660
rect 167644 4004 167696 4010
rect 167644 3946 167696 3952
rect 167748 3738 167776 70654
rect 167840 11830 167868 71810
rect 167932 14550 167960 71946
rect 168012 71936 168064 71942
rect 168012 71878 168064 71884
rect 168024 17474 168052 71878
rect 168116 22846 168144 72694
rect 168208 72690 168236 75140
rect 168300 73166 168328 75140
rect 168392 74934 168420 75140
rect 168380 74928 168432 74934
rect 168380 74870 168432 74876
rect 168484 74254 168512 75140
rect 168472 74248 168524 74254
rect 168472 74190 168524 74196
rect 168380 73296 168432 73302
rect 168380 73238 168432 73244
rect 168288 73160 168340 73166
rect 168288 73102 168340 73108
rect 168196 72684 168248 72690
rect 168196 72626 168248 72632
rect 168196 72412 168248 72418
rect 168196 72354 168248 72360
rect 168208 71482 168236 72354
rect 168286 72312 168342 72321
rect 168286 72247 168342 72256
rect 168300 71641 168328 72247
rect 168392 71777 168420 73238
rect 168472 72820 168524 72826
rect 168472 72762 168524 72768
rect 168378 71768 168434 71777
rect 168378 71703 168434 71712
rect 168286 71632 168342 71641
rect 168286 71567 168342 71576
rect 168208 71454 168328 71482
rect 168196 71120 168248 71126
rect 168196 71062 168248 71068
rect 168208 24274 168236 71062
rect 168300 36650 168328 71454
rect 168484 69222 168512 72762
rect 168576 72758 168604 75140
rect 168564 72752 168616 72758
rect 168564 72694 168616 72700
rect 168668 70145 168696 75140
rect 168760 72826 168788 75140
rect 168852 73302 168880 75140
rect 168840 73296 168892 73302
rect 168840 73238 168892 73244
rect 168944 73114 168972 75140
rect 168852 73086 168972 73114
rect 168748 72820 168800 72826
rect 168748 72762 168800 72768
rect 168852 70394 168880 73086
rect 169036 72978 169064 75140
rect 169128 73137 169156 75140
rect 169114 73128 169170 73137
rect 169114 73063 169170 73072
rect 169114 72992 169170 73001
rect 168932 72956 168984 72962
rect 169036 72950 169114 72978
rect 169114 72927 169170 72936
rect 168932 72898 168984 72904
rect 168760 70366 168880 70394
rect 168760 70281 168788 70366
rect 168746 70272 168802 70281
rect 168746 70207 168802 70216
rect 168654 70136 168710 70145
rect 168654 70071 168710 70080
rect 168472 69216 168524 69222
rect 168472 69158 168524 69164
rect 168380 65816 168432 65822
rect 168380 65758 168432 65764
rect 168288 36644 168340 36650
rect 168288 36586 168340 36592
rect 168196 24268 168248 24274
rect 168196 24210 168248 24216
rect 168104 22840 168156 22846
rect 168104 22782 168156 22788
rect 168012 17468 168064 17474
rect 168012 17410 168064 17416
rect 167920 14544 167972 14550
rect 167920 14486 167972 14492
rect 167828 11824 167880 11830
rect 167828 11766 167880 11772
rect 167736 3732 167788 3738
rect 167736 3674 167788 3680
rect 168392 480 168420 65758
rect 168944 64874 168972 72898
rect 169220 72865 169248 75140
rect 169206 72856 169262 72865
rect 169206 72791 169262 72800
rect 169116 72344 169168 72350
rect 169116 72286 169168 72292
rect 168944 64846 169064 64874
rect 169036 10402 169064 64846
rect 169128 19990 169156 72286
rect 169208 72208 169260 72214
rect 169208 72150 169260 72156
rect 169220 35290 169248 72150
rect 169312 69290 169340 75140
rect 169404 70378 169432 75140
rect 169496 74633 169524 75140
rect 169588 74866 169616 75140
rect 169576 74860 169628 74866
rect 169576 74802 169628 74808
rect 169482 74624 169538 74633
rect 169482 74559 169538 74568
rect 169680 73710 169708 75140
rect 169772 74866 169800 75140
rect 169760 74860 169812 74866
rect 169760 74802 169812 74808
rect 169864 74497 169892 75140
rect 169850 74488 169906 74497
rect 169850 74423 169906 74432
rect 169956 74322 169984 75140
rect 170048 74390 170076 75140
rect 170036 74384 170088 74390
rect 170036 74326 170088 74332
rect 169944 74316 169996 74322
rect 169944 74258 169996 74264
rect 170140 74118 170168 75140
rect 170128 74112 170180 74118
rect 170128 74054 170180 74060
rect 169668 73704 169720 73710
rect 169668 73646 169720 73652
rect 169392 70372 169444 70378
rect 169392 70314 169444 70320
rect 169576 69352 169628 69358
rect 169576 69294 169628 69300
rect 169300 69284 169352 69290
rect 169300 69226 169352 69232
rect 169208 35284 169260 35290
rect 169208 35226 169260 35232
rect 169116 19984 169168 19990
rect 169116 19926 169168 19932
rect 169024 10396 169076 10402
rect 169024 10338 169076 10344
rect 169588 480 169616 69294
rect 170232 45558 170260 75140
rect 170324 63034 170352 75140
rect 170416 74633 170444 75482
rect 170508 74866 170536 75618
rect 170496 74860 170548 74866
rect 170496 74802 170548 74808
rect 170402 74624 170458 74633
rect 170402 74559 170458 74568
rect 170600 73574 170628 75618
rect 170692 75585 170720 75618
rect 170678 75576 170734 75585
rect 170678 75511 170734 75520
rect 170678 75440 170734 75449
rect 170678 75375 170734 75384
rect 170692 75342 170720 75375
rect 170680 75336 170732 75342
rect 170680 75278 170732 75284
rect 172428 75268 172480 75274
rect 172428 75210 172480 75216
rect 170680 74996 170732 75002
rect 170680 74938 170732 74944
rect 170956 74996 171008 75002
rect 170956 74938 171008 74944
rect 170692 74866 170720 74938
rect 170680 74860 170732 74866
rect 170680 74802 170732 74808
rect 170588 73568 170640 73574
rect 170588 73510 170640 73516
rect 170968 73506 170996 74938
rect 172440 74934 172468 75210
rect 172428 74928 172480 74934
rect 172428 74870 172480 74876
rect 173162 74352 173218 74361
rect 173162 74287 173218 74296
rect 171784 74112 171836 74118
rect 171784 74054 171836 74060
rect 171796 73778 171824 74054
rect 171784 73772 171836 73778
rect 171784 73714 171836 73720
rect 172704 73636 172756 73642
rect 172704 73578 172756 73584
rect 170956 73500 171008 73506
rect 170956 73442 171008 73448
rect 172152 73024 172204 73030
rect 172336 73024 172388 73030
rect 172204 72972 172336 72978
rect 172152 72966 172388 72972
rect 172164 72950 172376 72966
rect 172716 72894 172744 73578
rect 172704 72888 172756 72894
rect 172704 72830 172756 72836
rect 170494 71904 170550 71913
rect 170494 71839 170550 71848
rect 170404 70848 170456 70854
rect 170404 70790 170456 70796
rect 170312 63028 170364 63034
rect 170312 62970 170364 62976
rect 170220 45552 170272 45558
rect 170220 45494 170272 45500
rect 170416 3874 170444 70790
rect 170404 3868 170456 3874
rect 170404 3810 170456 3816
rect 170508 3466 170536 71839
rect 171784 71732 171836 71738
rect 171784 71674 171836 71680
rect 171876 71732 171928 71738
rect 171876 71674 171928 71680
rect 171796 71126 171824 71674
rect 171784 71120 171836 71126
rect 171784 71062 171836 71068
rect 171888 70786 171916 71674
rect 171876 70780 171928 70786
rect 171876 70722 171928 70728
rect 170770 68640 170826 68649
rect 170770 68575 170826 68584
rect 170588 67176 170640 67182
rect 170588 67118 170640 67124
rect 170600 3534 170628 67118
rect 170588 3528 170640 3534
rect 170588 3470 170640 3476
rect 170496 3460 170548 3466
rect 170496 3402 170548 3408
rect 170784 480 170812 68575
rect 171966 62792 172022 62801
rect 171966 62727 172022 62736
rect 171980 480 172008 62727
rect 173176 480 173204 74287
rect 175292 73166 175320 76502
rect 175280 73160 175332 73166
rect 175280 73102 175332 73108
rect 173254 67144 173310 67153
rect 173254 67079 173310 67088
rect 173268 3602 173296 67079
rect 175462 64152 175518 64161
rect 175462 64087 175518 64096
rect 174266 52048 174322 52057
rect 174266 51983 174322 51992
rect 173256 3596 173308 3602
rect 173256 3538 173308 3544
rect 174280 480 174308 51983
rect 175476 480 175504 64087
rect 176660 58948 176712 58954
rect 176660 58890 176712 58896
rect 176672 480 176700 58890
rect 177040 33969 177068 132495
rect 177316 72690 177344 210394
rect 177868 121281 177896 214775
rect 188342 205728 188398 205737
rect 188342 205663 188398 205672
rect 185582 165880 185638 165889
rect 185582 165815 185638 165824
rect 178774 148336 178830 148345
rect 178774 148271 178830 148280
rect 178682 146976 178738 146985
rect 178682 146911 178738 146920
rect 178222 145616 178278 145625
rect 178222 145551 178278 145560
rect 178132 135924 178184 135930
rect 178132 135866 178184 135872
rect 178038 134328 178094 134337
rect 178038 134263 178094 134272
rect 178052 129713 178080 134263
rect 178038 129704 178094 129713
rect 178038 129639 178094 129648
rect 177854 121272 177910 121281
rect 177854 121207 177910 121216
rect 178144 110401 178172 135866
rect 178236 119785 178264 145551
rect 178314 144120 178370 144129
rect 178314 144055 178370 144064
rect 178222 119776 178278 119785
rect 178222 119711 178278 119720
rect 178222 118824 178278 118833
rect 178222 118759 178278 118768
rect 178130 110392 178186 110401
rect 178130 110327 178186 110336
rect 178236 109041 178264 118759
rect 178328 118289 178356 144055
rect 178406 142896 178462 142905
rect 178406 142831 178462 142840
rect 178314 118280 178370 118289
rect 178314 118215 178370 118224
rect 178420 116793 178448 142831
rect 178590 138680 178646 138689
rect 178590 138615 178646 138624
rect 178498 136232 178554 136241
rect 178498 136167 178554 136176
rect 178406 116784 178462 116793
rect 178406 116719 178462 116728
rect 178512 113121 178540 136167
rect 178604 115297 178632 138615
rect 178696 122505 178724 146911
rect 178788 124137 178816 148271
rect 178958 131200 179014 131209
rect 178958 131135 179014 131144
rect 178774 124128 178830 124137
rect 178774 124063 178830 124072
rect 178682 122496 178738 122505
rect 178682 122431 178738 122440
rect 178590 115288 178646 115297
rect 178590 115223 178646 115232
rect 178498 113112 178554 113121
rect 178498 113047 178554 113056
rect 178222 109032 178278 109041
rect 178222 108967 178278 108976
rect 177396 99408 177448 99414
rect 177396 99350 177448 99356
rect 177408 75682 177436 99350
rect 178498 86184 178554 86193
rect 178498 86119 178554 86128
rect 178512 80889 178540 86119
rect 178498 80880 178554 80889
rect 178498 80815 178554 80824
rect 178774 78704 178830 78713
rect 178774 78639 178830 78648
rect 177396 75676 177448 75682
rect 177396 75618 177448 75624
rect 178684 73092 178736 73098
rect 178684 73034 178736 73040
rect 178696 72962 178724 73034
rect 178684 72956 178736 72962
rect 178684 72898 178736 72904
rect 177304 72684 177356 72690
rect 177304 72626 177356 72632
rect 178684 64320 178736 64326
rect 178684 64262 178736 64268
rect 177856 56024 177908 56030
rect 177856 55966 177908 55972
rect 177026 33960 177082 33969
rect 177026 33895 177082 33904
rect 177868 480 177896 55966
rect 178696 3126 178724 64262
rect 178788 46345 178816 78639
rect 178866 76664 178922 76673
rect 178866 76599 178922 76608
rect 178880 64161 178908 76599
rect 178972 72321 179000 131135
rect 184202 126032 184258 126041
rect 184202 125967 184258 125976
rect 184216 82521 184244 125967
rect 185596 84017 185624 165815
rect 188356 85513 188384 205663
rect 207032 188358 207060 214540
rect 236012 214526 236578 214554
rect 266372 214526 266570 214554
rect 236012 189786 236040 214526
rect 266372 191146 266400 214526
rect 296732 213217 296760 214540
rect 296718 213208 296774 213217
rect 296718 213143 296774 213152
rect 266360 191140 266412 191146
rect 266360 191082 266412 191088
rect 236000 189780 236052 189786
rect 236000 189722 236052 189728
rect 207020 188352 207072 188358
rect 207020 188294 207072 188300
rect 327092 184249 327120 214540
rect 356532 212673 356560 214540
rect 386524 213217 386552 214540
rect 358082 213208 358138 213217
rect 358082 213143 358138 213152
rect 386510 213208 386566 213217
rect 386510 213143 386566 213152
rect 355322 212664 355378 212673
rect 355322 212599 355378 212608
rect 356518 212664 356574 212673
rect 356518 212599 356574 212608
rect 355336 186969 355364 212599
rect 355322 186960 355378 186969
rect 355322 186895 355378 186904
rect 327078 184240 327134 184249
rect 327078 184175 327134 184184
rect 358096 183569 358124 213143
rect 390572 212650 390600 214775
rect 390480 212622 390600 212650
rect 390480 211177 390508 212622
rect 387338 211168 387394 211177
rect 387338 211103 387394 211112
rect 390466 211168 390522 211177
rect 390466 211103 390522 211112
rect 387352 208457 387380 211103
rect 383658 208448 383714 208457
rect 383658 208383 383714 208392
rect 387338 208448 387394 208457
rect 387338 208383 387394 208392
rect 383672 207074 383700 208383
rect 383580 207046 383700 207074
rect 383580 204377 383608 207046
rect 378138 204368 378194 204377
rect 378138 204303 378194 204312
rect 383566 204368 383622 204377
rect 383566 204303 383622 204312
rect 378152 202994 378180 204303
rect 378060 202966 378180 202994
rect 378060 201385 378088 202966
rect 375378 201376 375434 201385
rect 375378 201311 375434 201320
rect 378046 201376 378102 201385
rect 378046 201311 378102 201320
rect 375392 198801 375420 201311
rect 375378 198792 375434 198801
rect 375378 198727 375434 198736
rect 369858 198656 369914 198665
rect 369858 198591 369914 198600
rect 369872 196058 369900 198591
rect 369780 196030 369900 196058
rect 369780 193905 369808 196030
rect 363602 193896 363658 193905
rect 363602 193831 363658 193840
rect 369766 193896 369822 193905
rect 369766 193831 369822 193840
rect 363616 186425 363644 193831
rect 360842 186416 360898 186425
rect 360842 186351 360898 186360
rect 363602 186416 363658 186425
rect 363602 186351 363658 186360
rect 358082 183560 358138 183569
rect 358082 183495 358138 183504
rect 199382 179208 199438 179217
rect 199382 179143 199438 179152
rect 199396 151065 199424 179143
rect 360856 173913 360884 186351
rect 359462 173904 359518 173913
rect 359462 173839 359518 173848
rect 360842 173904 360898 173913
rect 360842 173839 360898 173848
rect 199382 151056 199438 151065
rect 199382 150991 199438 151000
rect 359476 149161 359504 173839
rect 355690 149152 355746 149161
rect 355690 149087 355746 149096
rect 359462 149152 359518 149161
rect 359462 149087 359518 149096
rect 355704 142225 355732 149087
rect 351918 142216 351974 142225
rect 351918 142151 351974 142160
rect 355690 142216 355746 142225
rect 355690 142151 355746 142160
rect 351932 138145 351960 142151
rect 349158 138136 349214 138145
rect 349158 138071 349214 138080
rect 351918 138136 351974 138145
rect 351918 138071 351974 138080
rect 349172 136762 349200 138071
rect 349080 136734 349200 136762
rect 349080 135153 349108 136734
rect 345662 135144 345718 135153
rect 345662 135079 345718 135088
rect 349066 135144 349122 135153
rect 349066 135079 349122 135088
rect 345676 116521 345704 135079
rect 337382 116512 337438 116521
rect 337382 116447 337438 116456
rect 345662 116512 345718 116521
rect 345662 116447 345718 116456
rect 337396 109041 337424 116447
rect 331218 109032 331274 109041
rect 331218 108967 331274 108976
rect 337382 109032 337438 109041
rect 337382 108967 337438 108976
rect 331232 106865 331260 108967
rect 322938 106856 322994 106865
rect 322938 106791 322994 106800
rect 331218 106856 331274 106865
rect 331218 106791 331274 106800
rect 322952 106185 322980 106791
rect 322938 106176 322994 106185
rect 322938 106111 322994 106120
rect 396552 104825 396580 700431
rect 396630 700360 396686 700369
rect 396630 700295 396686 700304
rect 396644 214713 396672 700295
rect 396724 536852 396776 536858
rect 396724 536794 396776 536800
rect 396630 214704 396686 214713
rect 396630 214639 396686 214648
rect 396538 104816 396594 104825
rect 396538 104751 396594 104760
rect 188342 85504 188398 85513
rect 188342 85439 188398 85448
rect 185582 84008 185638 84017
rect 185582 83943 185638 83952
rect 184202 82512 184258 82521
rect 184202 82447 184258 82456
rect 228730 75304 228786 75313
rect 228730 75239 228786 75248
rect 196806 75168 196862 75177
rect 196806 75103 196862 75112
rect 179050 75032 179106 75041
rect 179050 74967 179106 74976
rect 178958 72312 179014 72321
rect 178958 72247 179014 72256
rect 178866 64152 178922 64161
rect 178866 64087 178922 64096
rect 178774 46336 178830 46345
rect 178774 46271 178830 46280
rect 178684 3120 178736 3126
rect 178684 3062 178736 3068
rect 179064 480 179092 74967
rect 194416 70916 194468 70922
rect 194416 70858 194468 70864
rect 189816 69624 189868 69630
rect 189816 69566 189868 69572
rect 181444 68808 181496 68814
rect 181444 68750 181496 68756
rect 180248 47864 180300 47870
rect 180248 47806 180300 47812
rect 180260 480 180288 47806
rect 181456 480 181484 68750
rect 184204 65748 184256 65754
rect 184204 65690 184256 65696
rect 183744 39568 183796 39574
rect 183744 39510 183796 39516
rect 182548 3120 182600 3126
rect 182548 3062 182600 3068
rect 182560 480 182588 3062
rect 183756 480 183784 39510
rect 184216 3398 184244 65690
rect 189722 61432 189778 61441
rect 189722 61367 189778 61376
rect 186136 53508 186188 53514
rect 186136 53450 186188 53456
rect 184940 49088 184992 49094
rect 184940 49030 184992 49036
rect 184204 3392 184256 3398
rect 184204 3334 184256 3340
rect 184952 480 184980 49030
rect 186148 480 186176 53450
rect 188528 46300 188580 46306
rect 188528 46242 188580 46248
rect 187332 3868 187384 3874
rect 187332 3810 187384 3816
rect 187344 480 187372 3810
rect 188540 480 188568 46242
rect 189736 480 189764 61367
rect 189828 3874 189856 69566
rect 192022 68504 192078 68513
rect 192022 68439 192078 68448
rect 190826 39400 190882 39409
rect 190826 39335 190882 39344
rect 189816 3868 189868 3874
rect 189816 3810 189868 3816
rect 190840 480 190868 39335
rect 192036 480 192064 68439
rect 193218 57488 193274 57497
rect 193218 57423 193274 57432
rect 193232 480 193260 57423
rect 194428 480 194456 70858
rect 195612 6044 195664 6050
rect 195612 5986 195664 5992
rect 195624 480 195652 5986
rect 196820 480 196848 75103
rect 214470 74896 214526 74905
rect 214470 74831 214526 74840
rect 208582 71224 208638 71233
rect 208582 71159 208638 71168
rect 200304 63096 200356 63102
rect 200304 63038 200356 63044
rect 197912 43648 197964 43654
rect 197912 43590 197964 43596
rect 197924 480 197952 43590
rect 199108 5160 199160 5166
rect 199108 5102 199160 5108
rect 199120 480 199148 5102
rect 200316 480 200344 63038
rect 207388 60240 207440 60246
rect 207388 60182 207440 60188
rect 201500 53440 201552 53446
rect 201500 53382 201552 53388
rect 201512 480 201540 53382
rect 203892 50652 203944 50658
rect 203892 50594 203944 50600
rect 202696 18828 202748 18834
rect 202696 18770 202748 18776
rect 202708 480 202736 18770
rect 203904 480 203932 50594
rect 206192 38140 206244 38146
rect 206192 38082 206244 38088
rect 205088 6112 205140 6118
rect 205088 6054 205140 6060
rect 205100 480 205128 6054
rect 206204 480 206232 38082
rect 207400 480 207428 60182
rect 208596 480 208624 71159
rect 213368 68740 213420 68746
rect 213368 68682 213420 68688
rect 210974 55992 211030 56001
rect 210974 55927 211030 55936
rect 209778 27024 209834 27033
rect 209778 26959 209834 26968
rect 209792 480 209820 26959
rect 210988 480 211016 55927
rect 212172 42288 212224 42294
rect 212172 42230 212224 42236
rect 212184 480 212212 42230
rect 213380 480 213408 68682
rect 214484 480 214512 74831
rect 218058 74760 218114 74769
rect 218058 74695 218114 74704
rect 216864 54800 216916 54806
rect 216864 54742 216916 54748
rect 215668 40928 215720 40934
rect 215668 40870 215720 40876
rect 215680 480 215708 40870
rect 216876 480 216904 54742
rect 218072 480 218100 74695
rect 227534 68368 227590 68377
rect 227534 68303 227590 68312
rect 221556 61532 221608 61538
rect 221556 61474 221608 61480
rect 219256 32700 219308 32706
rect 219256 32642 219308 32648
rect 219268 480 219296 32642
rect 220452 17536 220504 17542
rect 220452 17478 220504 17484
rect 220464 480 220492 17478
rect 221568 480 221596 61474
rect 225144 57452 225196 57458
rect 225144 57394 225196 57400
rect 223948 28620 224000 28626
rect 223948 28562 224000 28568
rect 222752 16176 222804 16182
rect 222752 16118 222804 16124
rect 222764 480 222792 16118
rect 223960 480 223988 28562
rect 225156 480 225184 57394
rect 226338 25664 226394 25673
rect 226338 25599 226394 25608
rect 226352 480 226380 25599
rect 227548 480 227576 68303
rect 228744 480 228772 75239
rect 235816 74860 235868 74866
rect 235816 74802 235868 74808
rect 232226 74216 232282 74225
rect 232226 74151 232282 74160
rect 231032 21684 231084 21690
rect 231032 21626 231084 21632
rect 229836 3392 229888 3398
rect 229836 3334 229888 3340
rect 229848 480 229876 3334
rect 231044 480 231072 21626
rect 232240 480 232268 74151
rect 234620 46232 234672 46238
rect 234620 46174 234672 46180
rect 233424 31340 233476 31346
rect 233424 31282 233476 31288
rect 233436 480 233464 31282
rect 234632 480 234660 46174
rect 235828 480 235856 74802
rect 249984 74792 250036 74798
rect 249984 74734 250036 74740
rect 247592 70984 247644 70990
rect 247592 70926 247644 70932
rect 241704 68672 241756 68678
rect 241704 68614 241756 68620
rect 239312 60172 239364 60178
rect 239312 60114 239364 60120
rect 237012 24472 237064 24478
rect 237012 24414 237064 24420
rect 237024 480 237052 24414
rect 238116 18760 238168 18766
rect 238116 18702 238168 18708
rect 238128 480 238156 18702
rect 239324 480 239352 60114
rect 240508 13388 240560 13394
rect 240508 13330 240560 13336
rect 240520 480 240548 13330
rect 241716 480 241744 68614
rect 242898 54632 242954 54641
rect 242898 54567 242954 54576
rect 242912 480 242940 54567
rect 246394 51912 246450 51921
rect 246394 51847 246450 51856
rect 244094 36680 244150 36689
rect 244094 36615 244150 36624
rect 244108 480 244136 36615
rect 245198 11928 245254 11937
rect 245198 11863 245254 11872
rect 245212 480 245240 11863
rect 246408 480 246436 51847
rect 247604 480 247632 70926
rect 248788 6860 248840 6866
rect 248788 6802 248840 6808
rect 248800 480 248828 6802
rect 249996 480 250024 74734
rect 285404 74724 285456 74730
rect 285404 74666 285456 74672
rect 267738 74080 267794 74089
rect 267738 74015 267794 74024
rect 251180 71664 251232 71670
rect 251180 71606 251232 71612
rect 251192 480 251220 71606
rect 253480 71596 253532 71602
rect 253480 71538 253532 71544
rect 252376 6792 252428 6798
rect 252376 6734 252428 6740
rect 252388 480 252416 6734
rect 253492 480 253520 71538
rect 262954 69728 263010 69737
rect 262954 69663 263010 69672
rect 259460 36712 259512 36718
rect 259460 36654 259512 36660
rect 254676 6724 254728 6730
rect 254676 6666 254728 6672
rect 254688 480 254716 6666
rect 258264 6656 258316 6662
rect 258264 6598 258316 6604
rect 255870 6488 255926 6497
rect 255870 6423 255926 6432
rect 255884 480 255912 6423
rect 257068 4140 257120 4146
rect 257068 4082 257120 4088
rect 257080 480 257108 4082
rect 258276 480 258304 6598
rect 259472 480 259500 36654
rect 261760 6588 261812 6594
rect 261760 6530 261812 6536
rect 260656 4072 260708 4078
rect 260656 4014 260708 4020
rect 260668 480 260696 4014
rect 261772 480 261800 6530
rect 262968 480 262996 69663
rect 266544 20256 266596 20262
rect 266544 20198 266596 20204
rect 265348 7812 265400 7818
rect 265348 7754 265400 7760
rect 264150 3768 264206 3777
rect 264150 3703 264206 3712
rect 264164 480 264192 3703
rect 265360 480 265388 7754
rect 266556 480 266584 20198
rect 267752 480 267780 74015
rect 283104 71528 283156 71534
rect 283104 71470 283156 71476
rect 279514 64288 279570 64297
rect 279514 64223 279570 64232
rect 277124 58880 277176 58886
rect 277124 58822 277176 58828
rect 271236 57384 271288 57390
rect 271236 57326 271288 57332
rect 270040 40860 270092 40866
rect 270040 40802 270092 40808
rect 268844 28552 268896 28558
rect 268844 28494 268896 28500
rect 268856 480 268884 28494
rect 270052 480 270080 40802
rect 271248 480 271276 57326
rect 274824 54732 274876 54738
rect 274824 54674 274876 54680
rect 272432 35420 272484 35426
rect 272432 35362 272484 35368
rect 272444 480 272472 35362
rect 273628 33924 273680 33930
rect 273628 33866 273680 33872
rect 273640 480 273668 33866
rect 274836 480 274864 54674
rect 276020 14748 276072 14754
rect 276020 14690 276072 14696
rect 276032 480 276060 14690
rect 277136 480 277164 58822
rect 278318 50416 278374 50425
rect 278318 50351 278374 50360
rect 278332 480 278360 50351
rect 279528 480 279556 64223
rect 281906 49056 281962 49065
rect 281906 48991 281962 49000
rect 280710 19952 280766 19961
rect 280710 19887 280766 19896
rect 280724 480 280752 19887
rect 281920 480 281948 48991
rect 283116 480 283144 71470
rect 284300 20188 284352 20194
rect 284300 20130 284352 20136
rect 284312 480 284340 20130
rect 285416 480 285444 74666
rect 320916 74656 320968 74662
rect 320916 74598 320968 74604
rect 306746 73400 306802 73409
rect 306746 73335 306802 73344
rect 288992 71460 289044 71466
rect 288992 71402 289044 71408
rect 286600 39500 286652 39506
rect 286600 39442 286652 39448
rect 286612 480 286640 39442
rect 287796 22908 287848 22914
rect 287796 22850 287848 22856
rect 287808 480 287836 22850
rect 289004 480 289032 71402
rect 298466 67008 298522 67017
rect 298466 66943 298522 66952
rect 291384 47796 291436 47802
rect 291384 47738 291436 47744
rect 290188 14680 290240 14686
rect 290188 14622 290240 14628
rect 290200 480 290228 14622
rect 291396 480 291424 47738
rect 293684 32632 293736 32638
rect 293684 32574 293736 32580
rect 292580 3936 292632 3942
rect 292580 3878 292632 3884
rect 292592 480 292620 3878
rect 293696 480 293724 32574
rect 294880 20120 294932 20126
rect 294880 20062 294932 20068
rect 294892 480 294920 20062
rect 297270 9072 297326 9081
rect 297270 9007 297326 9016
rect 296074 3632 296130 3641
rect 296074 3567 296130 3576
rect 296088 480 296116 3567
rect 297284 480 297312 9007
rect 298480 480 298508 66943
rect 300768 38072 300820 38078
rect 300768 38014 300820 38020
rect 299662 3496 299718 3505
rect 299662 3431 299718 3440
rect 299676 480 299704 3431
rect 300780 480 300808 38014
rect 304356 25764 304408 25770
rect 304356 25706 304408 25712
rect 301964 6520 302016 6526
rect 301964 6462 302016 6468
rect 301976 480 302004 6462
rect 303160 4004 303212 4010
rect 303160 3946 303212 3952
rect 303172 480 303200 3946
rect 304368 480 304396 25706
rect 305552 6452 305604 6458
rect 305552 6394 305604 6400
rect 305564 480 305592 6394
rect 306760 480 306788 73335
rect 307944 71392 307996 71398
rect 307944 71334 307996 71340
rect 307956 480 307984 71334
rect 311440 70236 311492 70242
rect 311440 70178 311492 70184
rect 310244 50584 310296 50590
rect 310244 50526 310296 50532
rect 309048 9308 309100 9314
rect 309048 9250 309100 9256
rect 309060 480 309088 9250
rect 310256 480 310284 50526
rect 311452 480 311480 70178
rect 317326 58712 317382 58721
rect 317326 58647 317382 58656
rect 313832 57316 313884 57322
rect 313832 57258 313884 57264
rect 312636 9240 312688 9246
rect 312636 9182 312688 9188
rect 312648 480 312676 9182
rect 313844 480 313872 57258
rect 315028 27124 315080 27130
rect 315028 27066 315080 27072
rect 315040 480 315068 27066
rect 316222 8936 316278 8945
rect 316222 8871 316278 8880
rect 316236 480 316264 8871
rect 317340 480 317368 58647
rect 319720 35352 319772 35358
rect 319720 35294 319772 35300
rect 318524 24404 318576 24410
rect 318524 24346 318576 24352
rect 318536 480 318564 24346
rect 319732 480 319760 35294
rect 320928 480 320956 74598
rect 343364 74588 343416 74594
rect 343364 74530 343416 74536
rect 332598 72720 332654 72729
rect 332598 72655 332654 72664
rect 332612 67114 332640 72655
rect 326804 67108 326856 67114
rect 326804 67050 326856 67056
rect 332600 67108 332652 67114
rect 332600 67050 332652 67056
rect 324412 54664 324464 54670
rect 324412 54606 324464 54612
rect 323308 16108 323360 16114
rect 323308 16050 323360 16056
rect 322112 5092 322164 5098
rect 322112 5034 322164 5040
rect 322124 480 322152 5034
rect 323320 480 323348 16050
rect 324424 480 324452 54606
rect 325608 13320 325660 13326
rect 325608 13262 325660 13268
rect 325620 480 325648 13262
rect 326816 480 326844 67050
rect 333886 66872 333942 66881
rect 333886 66807 333942 66816
rect 328000 51944 328052 51950
rect 328000 51886 328052 51892
rect 328012 480 328040 51886
rect 331586 47696 331642 47705
rect 331586 47631 331642 47640
rect 329196 10532 329248 10538
rect 329196 10474 329248 10480
rect 329208 480 329236 10474
rect 330392 5024 330444 5030
rect 330392 4966 330444 4972
rect 330404 480 330432 4966
rect 331600 480 331628 47631
rect 332690 22808 332746 22817
rect 332690 22743 332746 22752
rect 332704 480 332732 22743
rect 333900 480 333928 66807
rect 338672 60104 338724 60110
rect 338672 60046 338724 60052
rect 335082 46608 335138 46617
rect 335082 46543 335138 46552
rect 335096 480 335124 46543
rect 337476 32564 337528 32570
rect 337476 32506 337528 32512
rect 336280 14612 336332 14618
rect 336280 14554 336332 14560
rect 336292 480 336320 14554
rect 337488 480 337516 32506
rect 338684 480 338712 60046
rect 342168 53372 342220 53378
rect 342168 53314 342220 53320
rect 340972 21616 341024 21622
rect 340972 21558 341024 21564
rect 339868 7744 339920 7750
rect 339868 7686 339920 7692
rect 339880 480 339908 7686
rect 340984 480 341012 21558
rect 342180 480 342208 53314
rect 343376 480 343404 74530
rect 395342 73944 395398 73953
rect 395342 73879 395398 73888
rect 391848 71324 391900 71330
rect 391848 71266 391900 71272
rect 354036 70168 354088 70174
rect 354036 70110 354088 70116
rect 348056 67040 348108 67046
rect 348056 66982 348108 66988
rect 345756 49020 345808 49026
rect 345756 48962 345808 48968
rect 344560 21548 344612 21554
rect 344560 21490 344612 21496
rect 344572 480 344600 21490
rect 345768 480 345796 48962
rect 346952 3868 347004 3874
rect 346952 3810 347004 3816
rect 346964 480 346992 3810
rect 348068 480 348096 66982
rect 349250 44840 349306 44849
rect 349250 44775 349306 44784
rect 349264 480 349292 44775
rect 352838 43480 352894 43489
rect 352838 43415 352894 43424
rect 351642 21312 351698 21321
rect 351642 21247 351698 21256
rect 350446 10296 350502 10305
rect 350446 10231 350502 10240
rect 350460 480 350488 10231
rect 351656 480 351684 21247
rect 352852 480 352880 43415
rect 354048 480 354076 70110
rect 382372 70100 382424 70106
rect 382372 70042 382424 70048
rect 368202 69592 368258 69601
rect 368202 69527 368258 69536
rect 355232 66972 355284 66978
rect 355232 66914 355284 66920
rect 355244 480 355272 66914
rect 356336 62960 356388 62966
rect 356336 62902 356388 62908
rect 356348 480 356376 62902
rect 359924 55956 359976 55962
rect 359924 55898 359976 55904
rect 357532 31272 357584 31278
rect 357532 31214 357584 31220
rect 357544 480 357572 31214
rect 358728 21480 358780 21486
rect 358728 21422 358780 21428
rect 358740 480 358768 21422
rect 359936 480 359964 55898
rect 367008 50516 367060 50522
rect 367008 50458 367060 50464
rect 363512 47728 363564 47734
rect 363512 47670 363564 47676
rect 361120 42220 361172 42226
rect 361120 42162 361172 42168
rect 361132 480 361160 42162
rect 362316 38004 362368 38010
rect 362316 37946 362368 37952
rect 362328 480 362356 37946
rect 363524 480 363552 47670
rect 365812 21412 365864 21418
rect 365812 21354 365864 21360
rect 364616 9172 364668 9178
rect 364616 9114 364668 9120
rect 364628 480 364656 9114
rect 365824 480 365852 21354
rect 367020 480 367048 50458
rect 368216 480 368244 69527
rect 369400 66904 369452 66910
rect 369400 66846 369452 66852
rect 369412 480 369440 66846
rect 374092 61464 374144 61470
rect 374092 61406 374144 61412
rect 370594 40760 370650 40769
rect 370594 40695 370650 40704
rect 370608 480 370636 40695
rect 372896 28484 372948 28490
rect 372896 28426 372948 28432
rect 371700 25696 371752 25702
rect 371700 25638 371752 25644
rect 371712 480 371740 25638
rect 372908 480 372936 28426
rect 374104 480 374132 61406
rect 381176 60036 381228 60042
rect 381176 59978 381228 59984
rect 377680 51876 377732 51882
rect 377680 51818 377732 51824
rect 376484 18692 376536 18698
rect 376484 18634 376536 18640
rect 375288 16040 375340 16046
rect 375288 15982 375340 15988
rect 375300 480 375328 15982
rect 376496 480 376524 18634
rect 377692 480 377720 51818
rect 379980 27056 380032 27062
rect 379980 26998 380032 27004
rect 378876 15972 378928 15978
rect 378876 15914 378928 15920
rect 378888 480 378916 15914
rect 379992 480 380020 26998
rect 381188 480 381216 59978
rect 382384 480 382412 70042
rect 384762 46472 384818 46481
rect 384762 46407 384818 46416
rect 383568 20052 383620 20058
rect 383568 19994 383620 20000
rect 383580 480 383608 19994
rect 384776 480 384804 46407
rect 388258 39264 388314 39273
rect 388258 39199 388314 39208
rect 387154 33824 387210 33833
rect 387154 33759 387210 33768
rect 385958 11792 386014 11801
rect 385958 11727 386014 11736
rect 385972 480 386000 11727
rect 387168 480 387196 33759
rect 388272 480 388300 39199
rect 389456 24336 389508 24342
rect 389456 24278 389508 24284
rect 389468 480 389496 24278
rect 390652 4956 390704 4962
rect 390652 4898 390704 4904
rect 390664 480 390692 4898
rect 391860 480 391888 71266
rect 394240 62892 394292 62898
rect 394240 62834 394292 62840
rect 393044 15904 393096 15910
rect 393044 15846 393096 15852
rect 393056 480 393084 15846
rect 394252 480 394280 62834
rect 395356 480 395384 73879
rect 396736 72894 396764 536794
rect 397472 74254 397500 703520
rect 406382 700360 406438 700369
rect 397552 700324 397604 700330
rect 406382 700295 406438 700304
rect 397552 700266 397604 700272
rect 397460 74248 397512 74254
rect 397460 74190 397512 74196
rect 396724 72888 396776 72894
rect 396724 72830 396776 72836
rect 397564 72826 397592 700266
rect 405002 617536 405058 617545
rect 405002 617471 405058 617480
rect 403622 564360 403678 564369
rect 403622 564295 403678 564304
rect 400862 511320 400918 511329
rect 400862 511255 400918 511264
rect 399482 458144 399538 458153
rect 399482 458079 399538 458088
rect 399496 92449 399524 458079
rect 399574 219056 399630 219065
rect 399574 218991 399630 219000
rect 399588 203561 399616 218991
rect 399574 203552 399630 203561
rect 399574 203487 399630 203496
rect 400876 93809 400904 511255
rect 403636 95169 403664 564295
rect 405016 97889 405044 617471
rect 406396 100745 406424 700295
rect 413284 430636 413336 430642
rect 413284 430578 413336 430584
rect 411902 404968 411958 404977
rect 411902 404903 411958 404912
rect 409142 298752 409198 298761
rect 409142 298687 409198 298696
rect 407762 245576 407818 245585
rect 407762 245511 407818 245520
rect 406382 100736 406438 100745
rect 406382 100671 406438 100680
rect 405002 97880 405058 97889
rect 405002 97815 405058 97824
rect 403622 95160 403678 95169
rect 403622 95095 403678 95104
rect 400862 93800 400918 93809
rect 400862 93735 400918 93744
rect 399482 92440 399538 92449
rect 399482 92375 399538 92384
rect 407776 86873 407804 245511
rect 409156 88233 409184 298687
rect 410524 271924 410576 271930
rect 410524 271866 410576 271872
rect 409142 88224 409198 88233
rect 409142 88159 409198 88168
rect 407762 86864 407818 86873
rect 407762 86799 407818 86808
rect 410536 74458 410564 271866
rect 411916 91089 411944 404903
rect 411902 91080 411958 91089
rect 411902 91015 411958 91024
rect 413296 74526 413324 430578
rect 413664 136105 413692 703520
rect 429856 700641 429884 703520
rect 416042 700632 416098 700641
rect 416042 700567 416098 700576
rect 429842 700632 429898 700641
rect 429842 700567 429898 700576
rect 414662 700496 414718 700505
rect 414662 700431 414718 700440
rect 413650 136096 413706 136105
rect 413650 136031 413706 136040
rect 414676 102105 414704 700431
rect 416056 103465 416084 700567
rect 422944 590708 422996 590714
rect 422944 590650 422996 590656
rect 418804 484424 418856 484430
rect 418804 484366 418856 484372
rect 417424 324352 417476 324358
rect 417424 324294 417476 324300
rect 416042 103456 416098 103465
rect 416042 103391 416098 103400
rect 414662 102096 414718 102105
rect 414662 102031 414718 102040
rect 417436 75818 417464 324294
rect 417424 75812 417476 75818
rect 417424 75754 417476 75760
rect 413284 74520 413336 74526
rect 413284 74462 413336 74468
rect 410524 74452 410576 74458
rect 410524 74394 410576 74400
rect 418816 72962 418844 484366
rect 421564 378208 421616 378214
rect 421564 378150 421616 378156
rect 420182 351928 420238 351937
rect 420182 351863 420238 351872
rect 420196 89729 420224 351863
rect 420182 89720 420238 89729
rect 420182 89655 420238 89664
rect 421576 75886 421604 378150
rect 421564 75880 421616 75886
rect 421564 75822 421616 75828
rect 422956 73030 422984 590650
rect 446402 471472 446458 471481
rect 446402 471407 446458 471416
rect 442264 444440 442316 444446
rect 442264 444382 442316 444388
rect 439502 418296 439558 418305
rect 439502 418231 439558 418240
rect 433982 365120 434038 365129
rect 433982 365055 434038 365064
rect 429842 258904 429898 258913
rect 429842 258839 429898 258848
rect 429856 153785 429884 258839
rect 433996 156641 434024 365055
rect 438122 312080 438178 312089
rect 438122 312015 438178 312024
rect 433982 156632 434038 156641
rect 433982 156567 434038 156576
rect 438136 155281 438164 312015
rect 438122 155272 438178 155281
rect 438122 155207 438178 155216
rect 429842 153776 429898 153785
rect 429842 153711 429898 153720
rect 439516 142769 439544 418231
rect 442276 181393 442304 444382
rect 442262 181384 442318 181393
rect 442262 181319 442318 181328
rect 439502 142760 439558 142769
rect 439502 142695 439558 142704
rect 446416 137329 446444 471407
rect 446402 137320 446458 137329
rect 446402 137255 446458 137264
rect 462332 75274 462360 703520
rect 478524 195265 478552 703520
rect 494808 700505 494836 703520
rect 494794 700496 494850 700505
rect 494794 700431 494850 700440
rect 478510 195256 478566 195265
rect 478510 195191 478566 195200
rect 527192 76566 527220 703520
rect 543476 141409 543504 703520
rect 559668 700369 559696 703520
rect 559654 700360 559710 700369
rect 559654 700295 559710 700304
rect 580354 697232 580410 697241
rect 580354 697167 580410 697176
rect 544382 670712 544438 670721
rect 544382 670647 544438 670656
rect 543462 141400 543518 141409
rect 543462 141335 543518 141344
rect 544396 99385 544424 670647
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 579710 591016 579766 591025
rect 579710 590951 579766 590960
rect 579724 590714 579752 590951
rect 579712 590708 579764 590714
rect 579712 590650 579764 590656
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 580184 444446 580212 444751
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579632 324358 579660 325207
rect 579620 324352 579672 324358
rect 579620 324294 579672 324300
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579632 271930 579660 272167
rect 579620 271924 579672 271930
rect 579620 271866 579672 271872
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 544382 99376 544438 99385
rect 580172 99350 580224 99356
rect 544382 99311 544438 99320
rect 527180 76560 527232 76566
rect 527180 76502 527232 76508
rect 462320 75268 462372 75274
rect 462320 75210 462372 75216
rect 580276 75206 580304 643991
rect 580368 210458 580396 697167
rect 580538 683904 580594 683913
rect 580538 683839 580594 683848
rect 580446 630864 580502 630873
rect 580446 630799 580502 630808
rect 580356 210452 580408 210458
rect 580356 210394 580408 210400
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580264 75200 580316 75206
rect 580264 75142 580316 75148
rect 484032 74180 484084 74186
rect 484032 74122 484084 74128
rect 480534 73808 480590 73817
rect 480534 73743 480590 73752
rect 422944 73024 422996 73030
rect 422944 72966 422996 72972
rect 418804 72956 418856 72962
rect 418804 72898 418856 72904
rect 397552 72820 397604 72826
rect 397552 72762 397604 72768
rect 445024 72616 445076 72622
rect 445024 72558 445076 72564
rect 396540 70032 396592 70038
rect 396540 69974 396592 69980
rect 396552 480 396580 69974
rect 403624 69964 403676 69970
rect 403624 69906 403676 69912
rect 397736 64252 397788 64258
rect 397736 64194 397788 64200
rect 397748 480 397776 64194
rect 398932 45008 398984 45014
rect 398932 44950 398984 44956
rect 398944 480 398972 44950
rect 402520 42152 402572 42158
rect 402520 42094 402572 42100
rect 401324 22840 401376 22846
rect 401324 22782 401376 22788
rect 400128 4888 400180 4894
rect 400128 4830 400180 4836
rect 400140 480 400168 4830
rect 401336 480 401364 22782
rect 402532 480 402560 42094
rect 403636 480 403664 69906
rect 407212 69896 407264 69902
rect 407212 69838 407264 69844
rect 406014 37904 406070 37913
rect 406014 37839 406070 37848
rect 404818 25528 404874 25537
rect 404818 25463 404874 25472
rect 404832 480 404860 25463
rect 406028 480 406056 37839
rect 407224 480 407252 69838
rect 439134 59936 439190 59945
rect 439134 59871 439190 59880
rect 409604 58812 409656 58818
rect 409604 58754 409656 58760
rect 408408 24268 408460 24274
rect 408408 24210 408460 24216
rect 408420 480 408448 24210
rect 409616 480 409644 58754
rect 427268 54596 427320 54602
rect 427268 54538 427320 54544
rect 413100 53304 413152 53310
rect 413100 53246 413152 53252
rect 410800 13252 410852 13258
rect 410800 13194 410852 13200
rect 410812 480 410840 13194
rect 411904 9104 411956 9110
rect 411904 9046 411956 9052
rect 411916 480 411944 9046
rect 413112 480 413140 53246
rect 416688 47660 416740 47666
rect 416688 47602 416740 47608
rect 414296 14476 414348 14482
rect 414296 14418 414348 14424
rect 414308 480 414336 14418
rect 415492 11824 415544 11830
rect 415492 11766 415544 11772
rect 415504 480 415532 11766
rect 416700 480 416728 47602
rect 420182 40624 420238 40633
rect 420182 40559 420238 40568
rect 418986 7576 419042 7585
rect 418986 7511 419042 7520
rect 417884 6384 417936 6390
rect 417884 6326 417936 6332
rect 417896 480 417924 6326
rect 419000 480 419028 7511
rect 420196 480 420224 40559
rect 423770 36544 423826 36553
rect 423770 36479 423826 36488
rect 421378 22672 421434 22681
rect 421378 22607 421434 22616
rect 421392 480 421420 22607
rect 422576 14544 422628 14550
rect 422576 14486 422628 14492
rect 422588 480 422616 14486
rect 423784 480 423812 36479
rect 424968 33856 425020 33862
rect 424968 33798 425020 33804
rect 424980 480 425008 33798
rect 426164 13184 426216 13190
rect 426164 13126 426216 13132
rect 426176 480 426204 13126
rect 427280 480 427308 54538
rect 436744 51808 436796 51814
rect 436744 51750 436796 51756
rect 437938 51776 437994 51785
rect 430856 50448 430908 50454
rect 430856 50390 430908 50396
rect 429660 36644 429712 36650
rect 429660 36586 429712 36592
rect 428464 7676 428516 7682
rect 428464 7618 428516 7624
rect 428476 480 428504 7618
rect 429672 480 429700 36586
rect 430868 480 430896 50390
rect 434444 43580 434496 43586
rect 434444 43522 434496 43528
rect 432052 36576 432104 36582
rect 432052 36518 432104 36524
rect 432064 480 432092 36518
rect 433248 6316 433300 6322
rect 433248 6258 433300 6264
rect 433260 480 433288 6258
rect 434456 480 434484 43522
rect 435548 10464 435600 10470
rect 435548 10406 435600 10412
rect 435560 480 435588 10406
rect 436756 480 436784 51750
rect 437938 51711 437994 51720
rect 437952 480 437980 51711
rect 439148 480 439176 59871
rect 442632 47592 442684 47598
rect 442632 47534 442684 47540
rect 441526 35320 441582 35329
rect 441526 35255 441582 35264
rect 440330 30968 440386 30977
rect 440330 30903 440386 30912
rect 440344 480 440372 30903
rect 441540 480 441568 35255
rect 442644 480 442672 47534
rect 443828 17468 443880 17474
rect 443828 17410 443880 17416
rect 443840 480 443868 17410
rect 445036 480 445064 72558
rect 471244 72548 471296 72554
rect 471244 72490 471296 72496
rect 448612 71256 448664 71262
rect 448612 71198 448664 71204
rect 446220 65680 446272 65686
rect 446220 65622 446272 65628
rect 446232 480 446260 65622
rect 447416 44940 447468 44946
rect 447416 44882 447468 44888
rect 447428 480 447456 44882
rect 448624 480 448652 71198
rect 466276 69828 466328 69834
rect 466276 69770 466328 69776
rect 461584 68604 461636 68610
rect 461584 68546 461636 68552
rect 453304 61396 453356 61402
rect 453304 61338 453356 61344
rect 449808 28416 449860 28422
rect 449808 28358 449860 28364
rect 449820 480 449848 28358
rect 450912 19984 450964 19990
rect 450912 19926 450964 19932
rect 450924 480 450952 19926
rect 452108 3800 452160 3806
rect 452108 3742 452160 3748
rect 452120 480 452148 3742
rect 453316 480 453344 61338
rect 456890 35184 456946 35193
rect 456890 35119 456946 35128
rect 454500 29708 454552 29714
rect 454500 29650 454552 29656
rect 454512 480 454540 29650
rect 455696 3664 455748 3670
rect 455696 3606 455748 3612
rect 455708 480 455736 3606
rect 456904 480 456932 35119
rect 460388 29640 460440 29646
rect 460388 29582 460440 29588
rect 458088 10396 458140 10402
rect 458088 10338 458140 10344
rect 458100 480 458128 10338
rect 459190 3360 459246 3369
rect 459190 3295 459246 3304
rect 459204 480 459232 3295
rect 460400 480 460428 29582
rect 461596 480 461624 68546
rect 465172 35284 465224 35290
rect 465172 35226 465224 35232
rect 463976 17400 464028 17406
rect 463976 17342 464028 17348
rect 462780 3732 462832 3738
rect 462780 3674 462832 3680
rect 462792 480 462820 3674
rect 463988 480 464016 17342
rect 465184 480 465212 35226
rect 466288 480 466316 69770
rect 469864 69760 469916 69766
rect 469864 69702 469916 69708
rect 468668 54528 468720 54534
rect 468668 54470 468720 54476
rect 467472 17332 467524 17338
rect 467472 17274 467524 17280
rect 467484 480 467512 17274
rect 468680 480 468708 54470
rect 469876 480 469904 69702
rect 471060 17264 471112 17270
rect 471060 17206 471112 17212
rect 471072 480 471100 17206
rect 471256 8294 471284 72490
rect 475382 68232 475438 68241
rect 475382 68167 475438 68176
rect 472256 67108 472308 67114
rect 472256 67050 472308 67056
rect 471244 8288 471296 8294
rect 471244 8230 471296 8236
rect 472268 480 472296 67050
rect 472622 58576 472678 58585
rect 472622 58511 472678 58520
rect 472636 19825 472664 58511
rect 474554 57352 474610 57361
rect 474554 57287 474610 57296
rect 472622 19816 472678 19825
rect 472622 19751 472678 19760
rect 473450 6352 473506 6361
rect 473450 6287 473506 6296
rect 473464 480 473492 6287
rect 474568 480 474596 57287
rect 475396 3670 475424 68167
rect 478144 9036 478196 9042
rect 478144 8978 478196 8984
rect 476946 6216 477002 6225
rect 476946 6151 477002 6160
rect 475384 3664 475436 3670
rect 475384 3606 475436 3612
rect 475752 3596 475804 3602
rect 475752 3538 475804 3544
rect 475764 480 475792 3538
rect 476960 480 476988 6151
rect 478156 480 478184 8978
rect 479340 8288 479392 8294
rect 479340 8230 479392 8236
rect 479352 480 479380 8230
rect 480548 480 480576 73743
rect 481732 43512 481784 43518
rect 481732 43454 481784 43460
rect 481744 480 481772 43454
rect 482836 11756 482888 11762
rect 482836 11698 482888 11704
rect 482848 480 482876 11698
rect 484044 480 484072 74122
rect 515956 74112 516008 74118
rect 515956 74054 516008 74060
rect 505376 73228 505428 73234
rect 505376 73170 505428 73176
rect 501786 72584 501842 72593
rect 501786 72519 501842 72528
rect 497096 69692 497148 69698
rect 497096 69634 497148 69640
rect 487620 65612 487672 65618
rect 487620 65554 487672 65560
rect 486424 40792 486476 40798
rect 486424 40734 486476 40740
rect 485228 31204 485280 31210
rect 485228 31146 485280 31152
rect 485240 480 485268 31146
rect 486436 480 486464 40734
rect 487632 480 487660 65554
rect 491116 65544 491168 65550
rect 491116 65486 491168 65492
rect 488816 28348 488868 28354
rect 488816 28290 488868 28296
rect 488828 480 488856 28290
rect 489918 15872 489974 15881
rect 489918 15807 489974 15816
rect 489932 480 489960 15807
rect 491128 480 491156 65486
rect 494702 54496 494758 54505
rect 494702 54431 494758 54440
rect 492310 26888 492366 26897
rect 492310 26823 492366 26832
rect 492324 480 492352 26823
rect 493506 4856 493562 4865
rect 493506 4791 493562 4800
rect 493520 480 493548 4791
rect 494716 480 494744 54431
rect 495900 35216 495952 35222
rect 495900 35158 495952 35164
rect 495912 480 495940 35158
rect 497108 480 497136 69634
rect 500592 44872 500644 44878
rect 500592 44814 500644 44820
rect 499396 40724 499448 40730
rect 499396 40666 499448 40672
rect 498200 4820 498252 4826
rect 498200 4762 498252 4768
rect 498212 480 498240 4762
rect 499408 480 499436 40666
rect 500604 480 500632 44814
rect 501800 480 501828 72519
rect 504180 71188 504232 71194
rect 504180 71130 504232 71136
rect 502984 25628 503036 25634
rect 502984 25570 503036 25576
rect 502996 480 503024 25570
rect 504192 480 504220 71130
rect 505388 480 505416 73170
rect 512458 55856 512514 55865
rect 512458 55791 512514 55800
rect 508504 51740 508556 51746
rect 508504 51682 508556 51688
rect 506480 39432 506532 39438
rect 506480 39374 506532 39380
rect 506492 480 506520 39374
rect 507676 26988 507728 26994
rect 507676 26930 507728 26936
rect 507688 480 507716 26930
rect 508516 3602 508544 51682
rect 511262 50280 511318 50289
rect 511262 50215 511318 50224
rect 510068 24200 510120 24206
rect 510068 24142 510120 24148
rect 508504 3596 508556 3602
rect 508504 3538 508556 3544
rect 508872 3528 508924 3534
rect 508872 3470 508924 3476
rect 508884 480 508912 3470
rect 510080 480 510108 24142
rect 511276 480 511304 50215
rect 512472 480 512500 55791
rect 514760 43444 514812 43450
rect 514760 43386 514812 43392
rect 513564 22772 513616 22778
rect 513564 22714 513616 22720
rect 513576 480 513604 22714
rect 514772 480 514800 43386
rect 515968 480 515996 74054
rect 533712 74044 533764 74050
rect 533712 73986 533764 73992
rect 526626 65512 526682 65521
rect 526626 65447 526682 65456
rect 519544 64184 519596 64190
rect 519544 64126 519596 64132
rect 517152 33788 517204 33794
rect 517152 33730 517204 33736
rect 517164 480 517192 33730
rect 518348 32496 518400 32502
rect 518348 32438 518400 32444
rect 518360 480 518388 32438
rect 519556 480 519584 64126
rect 523040 62824 523092 62830
rect 523040 62766 523092 62772
rect 520740 32428 520792 32434
rect 520740 32370 520792 32376
rect 520752 480 520780 32370
rect 521844 25560 521896 25566
rect 521844 25502 521896 25508
rect 521856 480 521884 25502
rect 523052 480 523080 62766
rect 525432 42084 525484 42090
rect 525432 42026 525484 42032
rect 524236 3596 524288 3602
rect 524236 3538 524288 3544
rect 524248 480 524276 3538
rect 525444 480 525472 42026
rect 526640 480 526668 65447
rect 530122 57216 530178 57225
rect 530122 57151 530178 57160
rect 529018 14512 529074 14521
rect 529018 14447 529074 14456
rect 527822 11656 527878 11665
rect 527822 11591 527878 11600
rect 527836 480 527864 11591
rect 529032 480 529060 14447
rect 530136 480 530164 57151
rect 532516 24132 532568 24138
rect 532516 24074 532568 24080
rect 531320 8968 531372 8974
rect 531320 8910 531372 8916
rect 531332 480 531360 8910
rect 532528 480 532556 24074
rect 533724 480 533752 73986
rect 551468 73976 551520 73982
rect 551468 73918 551520 73924
rect 537208 73908 537260 73914
rect 537208 73850 537260 73856
rect 536104 31136 536156 31142
rect 536104 31078 536156 31084
rect 534908 10328 534960 10334
rect 534908 10270 534960 10276
rect 534920 480 534948 10270
rect 536116 480 536144 31078
rect 537220 480 537248 73850
rect 538404 71120 538456 71126
rect 538404 71062 538456 71068
rect 538416 480 538444 71062
rect 545488 71052 545540 71058
rect 545488 70994 545540 71000
rect 544384 58744 544436 58750
rect 544384 58686 544436 58692
rect 540796 57248 540848 57254
rect 540796 57190 540848 57196
rect 539600 53236 539652 53242
rect 539600 53178 539652 53184
rect 539612 480 539640 53178
rect 540808 480 540836 57190
rect 543188 39364 543240 39370
rect 543188 39306 543240 39312
rect 541992 7608 542044 7614
rect 541992 7550 542044 7556
rect 542004 480 542032 7550
rect 543200 480 543228 39306
rect 544396 480 544424 58686
rect 545500 480 545528 70994
rect 547878 42120 547934 42129
rect 547878 42055 547934 42064
rect 546684 3664 546736 3670
rect 546684 3606 546736 3612
rect 546696 480 546724 3606
rect 547892 480 547920 42055
rect 549076 31068 549128 31074
rect 549076 31010 549128 31016
rect 549088 480 549116 31010
rect 550272 13116 550324 13122
rect 550272 13058 550324 13064
rect 550284 480 550312 13058
rect 551480 480 551508 73918
rect 554964 73840 555016 73846
rect 554964 73782 555016 73788
rect 553768 68536 553820 68542
rect 553768 68478 553820 68484
rect 552664 53168 552716 53174
rect 552664 53110 552716 53116
rect 552676 480 552704 53110
rect 553780 480 553808 68478
rect 554976 480 555004 73782
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580184 72078 580212 72927
rect 580264 72480 580316 72486
rect 580264 72422 580316 72428
rect 580172 72072 580224 72078
rect 580172 72014 580224 72020
rect 577502 71904 577558 71913
rect 577502 71839 577558 71848
rect 559746 71088 559802 71097
rect 559746 71023 559802 71032
rect 558552 55888 558604 55894
rect 558552 55830 558604 55836
rect 556160 6248 556212 6254
rect 556160 6190 556212 6196
rect 556172 480 556200 6190
rect 557356 6180 557408 6186
rect 557356 6122 557408 6128
rect 557368 480 557396 6122
rect 558564 480 558592 55830
rect 559760 480 559788 71023
rect 560852 68468 560904 68474
rect 560852 68410 560904 68416
rect 560864 480 560892 68410
rect 568028 68400 568080 68406
rect 568028 68342 568080 68348
rect 562048 50380 562100 50386
rect 562048 50322 562100 50328
rect 562060 480 562088 50322
rect 565634 48920 565690 48929
rect 565634 48855 565690 48864
rect 563242 29608 563298 29617
rect 563242 29543 563298 29552
rect 563256 480 563284 29543
rect 564438 18728 564494 18737
rect 564438 18663 564494 18672
rect 564452 480 564480 18663
rect 565648 480 565676 48855
rect 566832 28280 566884 28286
rect 566832 28222 566884 28228
rect 566844 480 566872 28222
rect 568040 480 568068 68342
rect 575112 68332 575164 68338
rect 575112 68274 575164 68280
rect 572720 58676 572772 58682
rect 572720 58618 572772 58624
rect 569132 53100 569184 53106
rect 569132 53042 569184 53048
rect 569144 480 569172 53042
rect 570328 26920 570380 26926
rect 570328 26862 570380 26868
rect 570340 480 570368 26862
rect 571524 18624 571576 18630
rect 571524 18566 571576 18572
rect 571536 480 571564 18566
rect 572732 480 572760 58618
rect 573916 37936 573968 37942
rect 573916 37878 573968 37884
rect 573928 480 573956 37878
rect 575124 480 575152 68274
rect 576122 64152 576178 64161
rect 576122 64087 576178 64096
rect 576136 6633 576164 64087
rect 576306 47560 576362 47569
rect 576306 47495 576362 47504
rect 576122 6624 576178 6633
rect 576122 6559 576178 6568
rect 576320 480 576348 47495
rect 577410 13016 577466 13025
rect 577410 12951 577466 12960
rect 577424 480 577452 12951
rect 577516 3330 577544 71839
rect 580276 33153 580304 72422
rect 580368 71641 580396 192471
rect 580460 149705 580488 630799
rect 580552 209001 580580 683839
rect 580722 577688 580778 577697
rect 580722 577623 580778 577632
rect 580630 524512 580686 524521
rect 580630 524447 580686 524456
rect 580538 208992 580594 209001
rect 580538 208927 580594 208936
rect 580538 152688 580594 152697
rect 580538 152623 580594 152632
rect 580446 149696 580502 149705
rect 580446 149631 580502 149640
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580460 71738 580488 112775
rect 580448 71732 580500 71738
rect 580448 71674 580500 71680
rect 580354 71632 580410 71641
rect 580354 71567 580410 71576
rect 580552 71505 580580 152623
rect 580644 135969 580672 524447
rect 580736 214577 580764 577623
rect 580814 232384 580870 232393
rect 580814 232319 580870 232328
rect 580722 214568 580778 214577
rect 580722 214503 580778 214512
rect 580630 135960 580686 135969
rect 580630 135895 580686 135904
rect 580828 72146 580856 232319
rect 580816 72140 580868 72146
rect 580816 72082 580868 72088
rect 580538 71496 580594 71505
rect 580538 71431 580594 71440
rect 580998 46200 581054 46209
rect 580998 46135 581054 46144
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 578606 18592 578662 18601
rect 578606 18527 578662 18536
rect 577504 3324 577556 3330
rect 577504 3266 577556 3272
rect 578620 480 578648 18527
rect 581012 480 581040 46135
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 582196 3324 582248 3330
rect 582196 3266 582248 3272
rect 582208 480 582236 3266
rect 583404 480 583432 3402
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 658144 3478 658200
rect 3238 606056 3294 606112
rect 3330 553832 3386 553888
rect 2778 449540 2834 449576
rect 2778 449520 2780 449540
rect 2780 449520 2832 449540
rect 2832 449520 2834 449540
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 2778 345344 2834 345400
rect 3330 293120 3386 293176
rect 3330 241032 3386 241088
rect 3330 214920 3386 214976
rect 3330 210296 3386 210352
rect 3146 188808 3202 188864
rect 3330 162832 3386 162888
rect 3330 162016 3386 162072
rect 3330 136720 3386 136776
rect 3330 84632 3386 84688
rect 3698 566888 3754 566944
rect 3514 501744 3570 501800
rect 3422 73072 3478 73128
rect 3606 423544 3662 423600
rect 4802 514800 4858 514856
rect 3698 384240 3754 384296
rect 3698 267144 3754 267200
rect 3606 214784 3662 214840
rect 3698 211792 3754 211848
rect 3606 149776 3662 149832
rect 3606 133048 3662 133104
rect 3606 131144 3662 131200
rect 2778 6468 2780 6488
rect 2780 6468 2832 6488
rect 2832 6468 2834 6488
rect 2778 6432 2834 6468
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 33904 3478 33960
rect 3422 32408 3478 32464
rect 3698 128424 3754 128480
rect 3790 127064 3846 127120
rect 4986 462576 5042 462632
rect 4802 117136 4858 117192
rect 3790 97552 3846 97608
rect 4986 118632 5042 118688
rect 15842 684256 15898 684312
rect 11702 410488 11758 410544
rect 11702 119992 11758 120048
rect 14462 358400 14518 358456
rect 18602 632032 18658 632088
rect 22742 579944 22798 580000
rect 18602 138624 18658 138680
rect 15842 136176 15898 136232
rect 15842 134272 15898 134328
rect 14462 121352 14518 121408
rect 17958 133048 18014 133104
rect 17958 126928 18014 126984
rect 15842 110608 15898 110664
rect 22834 254088 22890 254144
rect 22742 142840 22798 142896
rect 22834 124072 22890 124128
rect 26882 671200 26938 671256
rect 25502 475632 25558 475688
rect 25594 384240 25650 384296
rect 25502 145560 25558 145616
rect 25594 115776 25650 115832
rect 29642 619112 29698 619168
rect 26974 371320 27030 371376
rect 26974 146920 27030 146976
rect 31022 527856 31078 527912
rect 29734 319232 29790 319288
rect 29734 148280 29790 148336
rect 31114 306176 31170 306232
rect 31022 144064 31078 144120
rect 45374 700576 45430 700632
rect 44914 700440 44970 700496
rect 40498 141480 40554 141536
rect 31114 122712 31170 122768
rect 29642 113056 29698 113112
rect 26882 111696 26938 111752
rect 24306 110336 24362 110392
rect 21362 74432 21418 74488
rect 8114 72936 8170 72992
rect 43442 72800 43498 72856
rect 25502 72528 25558 72584
rect 18234 71032 18290 71088
rect 3698 58520 3754 58576
rect 3606 19352 3662 19408
rect 21822 66816 21878 66872
rect 18602 51720 18658 51776
rect 34794 66952 34850 67008
rect 38382 53080 38438 53136
rect 37922 48864 37978 48920
rect 40774 50224 40830 50280
rect 44730 224168 44786 224224
rect 44730 216144 44786 216200
rect 45098 226072 45154 226128
rect 45098 108976 45154 109032
rect 45742 700304 45798 700360
rect 45374 107480 45430 107536
rect 44914 106120 44970 106176
rect 70950 281560 71006 281616
rect 69662 280064 69718 280120
rect 70950 280064 71006 280120
rect 67822 275984 67878 276040
rect 69662 275984 69718 276040
rect 45834 224848 45890 224904
rect 66534 270408 66590 270464
rect 67822 270408 67878 270464
rect 65522 264968 65578 265024
rect 66534 264968 66590 265024
rect 64142 248376 64198 248432
rect 65522 248376 65578 248432
rect 53838 231104 53894 231160
rect 64142 231104 64198 231160
rect 68926 226208 68982 226264
rect 53838 224984 53894 225040
rect 77942 334600 77998 334656
rect 76562 320864 76618 320920
rect 77942 320864 77998 320920
rect 75274 291080 75330 291136
rect 76562 291080 76618 291136
rect 73250 288496 73306 288552
rect 75274 288496 75330 288552
rect 73250 281560 73306 281616
rect 98918 236680 98974 236736
rect 95238 230424 95294 230480
rect 98918 230424 98974 230480
rect 89166 226072 89222 226128
rect 154118 700576 154174 700632
rect 167642 440816 167698 440872
rect 164882 427896 164938 427952
rect 167642 427896 167698 427952
rect 153842 356632 153898 356688
rect 164882 356632 164938 356688
rect 145838 342080 145894 342136
rect 153842 342080 153898 342136
rect 142802 338000 142858 338056
rect 145838 338000 145894 338056
rect 218978 700440 219034 700496
rect 220082 700440 220138 700496
rect 235170 700440 235226 700496
rect 283838 700304 283894 700360
rect 364982 700440 365038 700496
rect 396538 700440 396594 700496
rect 348790 700304 348846 700360
rect 300122 699896 300178 699952
rect 303158 699896 303214 699952
rect 303158 697448 303214 697504
rect 309782 697448 309838 697504
rect 309782 690104 309838 690160
rect 312542 690104 312598 690160
rect 312542 685752 312598 685808
rect 315302 685752 315358 685808
rect 213182 644544 213238 644600
rect 220082 644544 220138 644600
rect 207662 589872 207718 589928
rect 315302 663856 315358 663912
rect 317418 663856 317474 663912
rect 317418 658824 317474 658880
rect 337382 658824 337438 658880
rect 337382 646448 337438 646504
rect 345018 646448 345074 646504
rect 345018 639648 345074 639704
rect 348422 639648 348478 639704
rect 213182 589872 213238 589928
rect 204902 551928 204958 551984
rect 207662 551928 207718 551984
rect 348422 525816 348478 525872
rect 351182 525816 351238 525872
rect 197266 480800 197322 480856
rect 204902 480800 204958 480856
rect 184202 478080 184258 478136
rect 197266 478080 197322 478136
rect 178682 457408 178738 457464
rect 184202 457408 184258 457464
rect 178682 440816 178738 440872
rect 351182 351056 351238 351112
rect 376022 351056 376078 351112
rect 376022 339360 376078 339416
rect 378782 339360 378838 339416
rect 170310 334600 170366 334656
rect 378782 332424 378838 332480
rect 384578 332424 384634 332480
rect 384578 329024 384634 329080
rect 395342 329024 395398 329080
rect 139398 323584 139454 323640
rect 142802 323584 142858 323640
rect 129002 316648 129058 316704
rect 139398 316648 139454 316704
rect 126242 301552 126298 301608
rect 129002 301552 129058 301608
rect 120814 287680 120870 287736
rect 126242 287680 126298 287736
rect 395342 285640 395398 285696
rect 396446 285640 396502 285696
rect 117962 282240 118018 282296
rect 120814 282240 120870 282296
rect 113822 272176 113878 272232
rect 117962 272176 118018 272232
rect 108302 266328 108358 266384
rect 113822 266328 113878 266384
rect 105542 253952 105598 254008
rect 108302 253952 108358 254008
rect 105542 236680 105598 236736
rect 105450 226208 105506 226264
rect 95238 224168 95294 224224
rect 46846 216144 46902 216200
rect 45834 215872 45890 215928
rect 46846 210432 46902 210488
rect 56598 210432 56654 210488
rect 56598 205672 56654 205728
rect 46202 201864 46258 201920
rect 149058 215872 149114 215928
rect 114374 214648 114430 214704
rect 58622 205672 58678 205728
rect 57886 193840 57942 193896
rect 58622 191664 58678 191720
rect 60002 191664 60058 191720
rect 60002 186360 60058 186416
rect 61382 186360 61438 186416
rect 88246 182008 88302 182064
rect 61382 167048 61438 167104
rect 62762 167048 62818 167104
rect 62762 144200 62818 144256
rect 70766 144200 70822 144256
rect 70766 140800 70822 140856
rect 73158 140800 73214 140856
rect 73158 134408 73214 134464
rect 46202 125432 46258 125488
rect 45742 104760 45798 104816
rect 44822 70216 44878 70272
rect 52550 64096 52606 64152
rect 53746 46144 53802 46200
rect 70306 58656 70362 58712
rect 72606 68176 72662 68232
rect 73802 50360 73858 50416
rect 74998 49000 75054 49056
rect 113730 137264 113786 137320
rect 114006 156576 114062 156632
rect 113914 142704 113970 142760
rect 113822 133184 113878 133240
rect 113822 129784 113878 129840
rect 113730 91024 113786 91080
rect 113914 89664 113970 89720
rect 114098 155216 114154 155272
rect 114006 88168 114062 88224
rect 114190 153720 114246 153776
rect 114098 86808 114154 86864
rect 114282 151000 114338 151056
rect 114190 85312 114246 85368
rect 115846 214512 115902 214568
rect 115754 208936 115810 208992
rect 114466 203496 114522 203552
rect 114374 103128 114430 103184
rect 114282 82320 114338 82376
rect 113822 80824 113878 80880
rect 115662 149640 115718 149696
rect 115478 141344 115534 141400
rect 115386 136040 115442 136096
rect 115386 101768 115442 101824
rect 115570 135904 115626 135960
rect 115478 98776 115534 98832
rect 115754 96668 115810 96724
rect 115662 95172 115718 95228
rect 116766 195200 116822 195256
rect 116490 129820 116492 129840
rect 116492 129820 116544 129840
rect 116544 129820 116546 129840
rect 116490 129784 116546 129820
rect 116490 100308 116492 100328
rect 116492 100308 116544 100328
rect 116544 100308 116546 100328
rect 116490 100272 116546 100308
rect 115846 93676 115902 93732
rect 115570 92384 115626 92440
rect 114466 83680 114522 83736
rect 114374 76608 114430 76664
rect 105726 71168 105782 71224
rect 104162 70080 104218 70136
rect 90362 69672 90418 69728
rect 87970 61376 88026 61432
rect 89166 6160 89222 6216
rect 91558 55800 91614 55856
rect 116490 78104 116546 78160
rect 116490 75520 116546 75576
rect 114466 75112 114522 75168
rect 114374 59608 114430 59664
rect 114466 58520 114522 58576
rect 116674 139304 116730 139360
rect 177854 214784 177910 214840
rect 390558 214784 390614 214840
rect 396446 214784 396502 214840
rect 149058 213152 149114 213208
rect 159362 213152 159418 213208
rect 162122 213152 162178 213208
rect 159362 209072 159418 209128
rect 143446 207032 143502 207088
rect 146298 207032 146354 207088
rect 134522 193840 134578 193896
rect 157246 186904 157302 186960
rect 152738 184184 152794 184240
rect 155958 183504 156014 183560
rect 154302 183368 154358 183424
rect 157246 183368 157302 183424
rect 133234 182028 133290 182064
rect 133234 182008 133236 182028
rect 133236 182008 133288 182028
rect 133288 182008 133290 182028
rect 136638 182028 136694 182064
rect 136638 182008 136640 182028
rect 136640 182008 136692 182028
rect 136692 182008 136694 182028
rect 117226 180648 117282 180704
rect 133234 180648 133290 180704
rect 136362 179460 136364 179480
rect 136364 179460 136416 179480
rect 136416 179460 136418 179480
rect 136362 179424 136418 179460
rect 138570 181328 138626 181384
rect 137834 181192 137890 181248
rect 138018 181076 138074 181112
rect 138754 181192 138810 181248
rect 138018 181056 138020 181076
rect 138020 181056 138072 181076
rect 138072 181056 138074 181076
rect 154486 181328 154542 181384
rect 140962 179696 141018 179752
rect 149886 179968 149942 180024
rect 146022 179560 146078 179616
rect 146298 179424 146354 179480
rect 151726 179832 151782 179888
rect 150990 179696 151046 179752
rect 176842 211792 176898 211848
rect 167642 209072 167698 209128
rect 167642 198736 167698 198792
rect 173162 198736 173218 198792
rect 173162 186360 173218 186416
rect 175278 210296 175334 210352
rect 155774 181736 155830 181792
rect 162122 181736 162178 181792
rect 155406 181328 155462 181384
rect 163042 181328 163098 181384
rect 155406 179968 155462 180024
rect 155498 179832 155554 179888
rect 155774 179696 155830 179752
rect 162766 179424 162822 179480
rect 142618 176024 142674 176080
rect 141882 172488 141938 172544
rect 139490 165144 139546 165200
rect 136086 162016 136142 162072
rect 136362 162016 136418 162072
rect 122470 137400 122526 137456
rect 125598 137536 125654 137592
rect 160466 161492 160522 161528
rect 160466 161472 160468 161492
rect 160468 161472 160520 161492
rect 160520 161472 160522 161492
rect 163226 161472 163282 161528
rect 139490 161064 139546 161120
rect 161570 152360 161626 152416
rect 163686 160656 163742 160712
rect 168378 162152 168434 162208
rect 167826 137400 167882 137456
rect 175922 186360 175978 186416
rect 175370 126928 175426 126984
rect 176750 162016 176806 162072
rect 176658 134408 176714 134464
rect 175922 118768 175978 118824
rect 176750 128288 176806 128344
rect 176934 141480 176990 141536
rect 176842 125432 176898 125488
rect 177026 132504 177082 132560
rect 176934 111696 176990 111752
rect 176658 107480 176714 107536
rect 117870 73072 117926 73128
rect 117870 72528 117926 72584
rect 116858 71984 116914 72040
rect 116674 69536 116730 69592
rect 117962 70352 118018 70408
rect 120262 72936 120318 72992
rect 120262 72664 120318 72720
rect 120078 71712 120134 71768
rect 121642 72664 121698 72720
rect 121458 70488 121514 70544
rect 121918 72936 121974 72992
rect 122378 71984 122434 72040
rect 122838 72392 122894 72448
rect 123206 72664 123262 72720
rect 123390 72528 123446 72584
rect 123666 73480 123722 73536
rect 123574 72800 123630 72856
rect 123758 72528 123814 72584
rect 123666 71032 123722 71088
rect 124310 73072 124366 73128
rect 124218 72664 124274 72720
rect 124586 72800 124642 72856
rect 124494 72664 124550 72720
rect 124402 72528 124458 72584
rect 125690 72800 125746 72856
rect 125598 72664 125654 72720
rect 126426 72528 126482 72584
rect 126702 72936 126758 72992
rect 126978 72800 127034 72856
rect 127254 72664 127310 72720
rect 127162 72528 127218 72584
rect 127346 72392 127402 72448
rect 128358 72800 128414 72856
rect 128450 72528 128506 72584
rect 128634 72664 128690 72720
rect 128542 69672 128598 69728
rect 129738 73072 129794 73128
rect 129830 72664 129886 72720
rect 129830 71168 129886 71224
rect 132406 72800 132462 72856
rect 132314 72664 132370 72720
rect 133694 72800 133750 72856
rect 133602 72664 133658 72720
rect 133510 72528 133566 72584
rect 133786 72392 133842 72448
rect 134062 72936 134118 72992
rect 134982 74296 135038 74352
rect 135074 72800 135130 72856
rect 134890 72664 134946 72720
rect 134798 72392 134854 72448
rect 135166 72528 135222 72584
rect 135442 74840 135498 74896
rect 136454 72800 136510 72856
rect 136362 72664 136418 72720
rect 136546 72528 136602 72584
rect 136270 72392 136326 72448
rect 136822 72256 136878 72312
rect 136270 48184 136326 48240
rect 137926 72800 137982 72856
rect 137834 72664 137890 72720
rect 137742 71440 137798 71496
rect 138202 71848 138258 71904
rect 138478 72120 138534 72176
rect 139122 73480 139178 73536
rect 139214 73344 139270 73400
rect 139306 73072 139362 73128
rect 139582 74160 139638 74216
rect 139582 72392 139638 72448
rect 139858 73208 139914 73264
rect 140502 73480 140558 73536
rect 140686 73616 140742 73672
rect 140410 73344 140466 73400
rect 140594 73344 140650 73400
rect 140042 17176 140098 17232
rect 138846 3304 138902 3360
rect 142066 73480 142122 73536
rect 142066 72256 142122 72312
rect 141974 69672 142030 69728
rect 142342 74024 142398 74080
rect 143354 72936 143410 72992
rect 143262 72800 143318 72856
rect 143170 72664 143226 72720
rect 143446 72528 143502 72584
rect 143722 72256 143778 72312
rect 144826 72800 144882 72856
rect 144734 72664 144790 72720
rect 144642 72528 144698 72584
rect 144826 72528 144882 72584
rect 144550 72392 144606 72448
rect 144826 72120 144882 72176
rect 145378 72936 145434 72992
rect 146206 72800 146262 72856
rect 146114 72664 146170 72720
rect 147310 72664 147366 72720
rect 147402 72120 147458 72176
rect 147494 71440 147550 71496
rect 147586 71304 147642 71360
rect 147770 72936 147826 72992
rect 147770 72120 147826 72176
rect 148690 73072 148746 73128
rect 148874 72800 148930 72856
rect 148782 72664 148838 72720
rect 148966 72528 149022 72584
rect 149242 65320 149298 65376
rect 149978 65592 150034 65648
rect 150162 72800 150218 72856
rect 150438 73072 150494 73128
rect 150346 72664 150402 72720
rect 151082 72392 151138 72448
rect 151082 71848 151138 71904
rect 151634 73888 151690 73944
rect 151542 72664 151598 72720
rect 151450 72528 151506 72584
rect 151726 72392 151782 72448
rect 152278 74568 152334 74624
rect 152738 72800 152794 72856
rect 151174 15816 151230 15872
rect 153106 73480 153162 73536
rect 153106 72936 153162 72992
rect 153014 72664 153070 72720
rect 153290 72936 153346 72992
rect 153842 72256 153898 72312
rect 154210 72800 154266 72856
rect 154302 72664 154358 72720
rect 154118 72392 154174 72448
rect 154486 72528 154542 72584
rect 155590 72800 155646 72856
rect 155774 72664 155830 72720
rect 155682 72528 155738 72584
rect 155866 72392 155922 72448
rect 156142 72276 156198 72312
rect 156142 72256 156144 72276
rect 156144 72256 156196 72276
rect 156196 72256 156198 72276
rect 155222 37984 155278 38040
rect 157246 72528 157302 72584
rect 156602 42064 156658 42120
rect 157154 71848 157210 71904
rect 157522 73072 157578 73128
rect 157706 74840 157762 74896
rect 157706 73208 157762 73264
rect 157982 73072 158038 73128
rect 157982 72664 158038 72720
rect 157982 72120 158038 72176
rect 158350 72664 158406 72720
rect 158534 72664 158590 72720
rect 158626 72528 158682 72584
rect 158442 72392 158498 72448
rect 158626 72392 158682 72448
rect 158350 72120 158406 72176
rect 158902 73752 158958 73808
rect 158902 73364 158958 73400
rect 158902 73344 158904 73364
rect 158904 73344 158956 73364
rect 158956 73344 158958 73364
rect 159178 72664 159234 72720
rect 159638 72664 159694 72720
rect 159914 72664 159970 72720
rect 159822 72528 159878 72584
rect 160282 72664 160338 72720
rect 160558 72392 160614 72448
rect 161202 73480 161258 73536
rect 161294 73208 161350 73264
rect 161018 72664 161074 72720
rect 160742 71304 160798 71360
rect 161386 72528 161442 72584
rect 162214 70352 162270 70408
rect 162582 73072 162638 73128
rect 162674 72664 162730 72720
rect 162490 72528 162546 72584
rect 162766 72392 162822 72448
rect 162766 70352 162822 70408
rect 163318 71848 163374 71904
rect 161294 3848 161350 3904
rect 163962 72528 164018 72584
rect 164146 72664 164202 72720
rect 164146 72528 164202 72584
rect 164054 72392 164110 72448
rect 165066 71032 165122 71088
rect 165342 72664 165398 72720
rect 165434 72528 165490 72584
rect 165526 72392 165582 72448
rect 165710 72528 165766 72584
rect 165710 72120 165766 72176
rect 165710 71848 165766 71904
rect 166538 72528 166594 72584
rect 166446 72392 166502 72448
rect 166354 72120 166410 72176
rect 166630 72120 166686 72176
rect 166814 73480 166870 73536
rect 166722 71984 166778 72040
rect 167550 74568 167606 74624
rect 167274 71440 167330 71496
rect 167182 71304 167238 71360
rect 168286 72256 168342 72312
rect 168378 71712 168434 71768
rect 168286 71576 168342 71632
rect 169114 73072 169170 73128
rect 169114 72936 169170 72992
rect 168746 70216 168802 70272
rect 168654 70080 168710 70136
rect 169206 72800 169262 72856
rect 169482 74568 169538 74624
rect 169850 74432 169906 74488
rect 170402 74568 170458 74624
rect 170678 75520 170734 75576
rect 170678 75384 170734 75440
rect 173162 74296 173218 74352
rect 170494 71848 170550 71904
rect 170770 68584 170826 68640
rect 171966 62736 172022 62792
rect 173254 67088 173310 67144
rect 175462 64096 175518 64152
rect 174266 51992 174322 52048
rect 188342 205672 188398 205728
rect 185582 165824 185638 165880
rect 178774 148280 178830 148336
rect 178682 146920 178738 146976
rect 178222 145560 178278 145616
rect 178038 134272 178094 134328
rect 178038 129648 178094 129704
rect 177854 121216 177910 121272
rect 178314 144064 178370 144120
rect 178222 119720 178278 119776
rect 178222 118768 178278 118824
rect 178130 110336 178186 110392
rect 178406 142840 178462 142896
rect 178314 118224 178370 118280
rect 178590 138624 178646 138680
rect 178498 136176 178554 136232
rect 178406 116728 178462 116784
rect 178958 131144 179014 131200
rect 178774 124072 178830 124128
rect 178682 122440 178738 122496
rect 178590 115232 178646 115288
rect 178498 113056 178554 113112
rect 178222 108976 178278 109032
rect 178498 86128 178554 86184
rect 178498 80824 178554 80880
rect 178774 78648 178830 78704
rect 177026 33904 177082 33960
rect 178866 76608 178922 76664
rect 184202 125976 184258 126032
rect 296718 213152 296774 213208
rect 358082 213152 358138 213208
rect 386510 213152 386566 213208
rect 355322 212608 355378 212664
rect 356518 212608 356574 212664
rect 355322 186904 355378 186960
rect 327078 184184 327134 184240
rect 387338 211112 387394 211168
rect 390466 211112 390522 211168
rect 383658 208392 383714 208448
rect 387338 208392 387394 208448
rect 378138 204312 378194 204368
rect 383566 204312 383622 204368
rect 375378 201320 375434 201376
rect 378046 201320 378102 201376
rect 375378 198736 375434 198792
rect 369858 198600 369914 198656
rect 363602 193840 363658 193896
rect 369766 193840 369822 193896
rect 360842 186360 360898 186416
rect 363602 186360 363658 186416
rect 358082 183504 358138 183560
rect 199382 179152 199438 179208
rect 359462 173848 359518 173904
rect 360842 173848 360898 173904
rect 199382 151000 199438 151056
rect 355690 149096 355746 149152
rect 359462 149096 359518 149152
rect 351918 142160 351974 142216
rect 355690 142160 355746 142216
rect 349158 138080 349214 138136
rect 351918 138080 351974 138136
rect 345662 135088 345718 135144
rect 349066 135088 349122 135144
rect 337382 116456 337438 116512
rect 345662 116456 345718 116512
rect 331218 108976 331274 109032
rect 337382 108976 337438 109032
rect 322938 106800 322994 106856
rect 331218 106800 331274 106856
rect 322938 106120 322994 106176
rect 396630 700304 396686 700360
rect 396630 214648 396686 214704
rect 396538 104760 396594 104816
rect 188342 85448 188398 85504
rect 185582 83952 185638 84008
rect 184202 82456 184258 82512
rect 228730 75248 228786 75304
rect 196806 75112 196862 75168
rect 179050 74976 179106 75032
rect 178958 72256 179014 72312
rect 178866 64096 178922 64152
rect 178774 46280 178830 46336
rect 189722 61376 189778 61432
rect 192022 68448 192078 68504
rect 190826 39344 190882 39400
rect 193218 57432 193274 57488
rect 214470 74840 214526 74896
rect 208582 71168 208638 71224
rect 210974 55936 211030 55992
rect 209778 26968 209834 27024
rect 218058 74704 218114 74760
rect 227534 68312 227590 68368
rect 226338 25608 226394 25664
rect 232226 74160 232282 74216
rect 242898 54576 242954 54632
rect 246394 51856 246450 51912
rect 244094 36624 244150 36680
rect 245198 11872 245254 11928
rect 267738 74024 267794 74080
rect 262954 69672 263010 69728
rect 255870 6432 255926 6488
rect 264150 3712 264206 3768
rect 279514 64232 279570 64288
rect 278318 50360 278374 50416
rect 281906 49000 281962 49056
rect 280710 19896 280766 19952
rect 306746 73344 306802 73400
rect 298466 66952 298522 67008
rect 297270 9016 297326 9072
rect 296074 3576 296130 3632
rect 299662 3440 299718 3496
rect 317326 58656 317382 58712
rect 316222 8880 316278 8936
rect 332598 72664 332654 72720
rect 333886 66816 333942 66872
rect 331586 47640 331642 47696
rect 332690 22752 332746 22808
rect 335082 46552 335138 46608
rect 395342 73888 395398 73944
rect 349250 44784 349306 44840
rect 352838 43424 352894 43480
rect 351642 21256 351698 21312
rect 350446 10240 350502 10296
rect 368202 69536 368258 69592
rect 370594 40704 370650 40760
rect 384762 46416 384818 46472
rect 388258 39208 388314 39264
rect 387154 33768 387210 33824
rect 385958 11736 386014 11792
rect 406382 700304 406438 700360
rect 405002 617480 405058 617536
rect 403622 564304 403678 564360
rect 400862 511264 400918 511320
rect 399482 458088 399538 458144
rect 399574 219000 399630 219056
rect 399574 203496 399630 203552
rect 411902 404912 411958 404968
rect 409142 298696 409198 298752
rect 407762 245520 407818 245576
rect 406382 100680 406438 100736
rect 405002 97824 405058 97880
rect 403622 95104 403678 95160
rect 400862 93744 400918 93800
rect 399482 92384 399538 92440
rect 409142 88168 409198 88224
rect 407762 86808 407818 86864
rect 411902 91024 411958 91080
rect 416042 700576 416098 700632
rect 429842 700576 429898 700632
rect 414662 700440 414718 700496
rect 413650 136040 413706 136096
rect 416042 103400 416098 103456
rect 414662 102040 414718 102096
rect 420182 351872 420238 351928
rect 420182 89664 420238 89720
rect 446402 471416 446458 471472
rect 439502 418240 439558 418296
rect 433982 365064 434038 365120
rect 429842 258848 429898 258904
rect 438122 312024 438178 312080
rect 433982 156576 434038 156632
rect 438122 155216 438178 155272
rect 429842 153720 429898 153776
rect 442262 181328 442318 181384
rect 439502 142704 439558 142760
rect 446402 137264 446458 137320
rect 494794 700440 494850 700496
rect 478510 195200 478566 195256
rect 559654 700304 559710 700360
rect 580354 697176 580410 697232
rect 544382 670656 544438 670712
rect 543462 141344 543518 141400
rect 580262 644000 580318 644056
rect 579710 590960 579766 591016
rect 580170 537784 580226 537840
rect 580170 484608 580226 484664
rect 580170 444760 580226 444816
rect 580170 431568 580226 431624
rect 580170 378392 580226 378448
rect 579618 325216 579674 325272
rect 579618 272176 579674 272232
rect 580170 99456 580226 99512
rect 544382 99320 544438 99376
rect 580538 683848 580594 683904
rect 580446 630808 580502 630864
rect 580354 192480 580410 192536
rect 480534 73752 480590 73808
rect 406014 37848 406070 37904
rect 404818 25472 404874 25528
rect 439134 59880 439190 59936
rect 420182 40568 420238 40624
rect 418986 7520 419042 7576
rect 423770 36488 423826 36544
rect 421378 22616 421434 22672
rect 437938 51720 437994 51776
rect 441526 35264 441582 35320
rect 440330 30912 440386 30968
rect 456890 35128 456946 35184
rect 459190 3304 459246 3360
rect 475382 68176 475438 68232
rect 472622 58520 472678 58576
rect 474554 57296 474610 57352
rect 472622 19760 472678 19816
rect 473450 6296 473506 6352
rect 476946 6160 477002 6216
rect 501786 72528 501842 72584
rect 489918 15816 489974 15872
rect 494702 54440 494758 54496
rect 492310 26832 492366 26888
rect 493506 4800 493562 4856
rect 512458 55800 512514 55856
rect 511262 50224 511318 50280
rect 526626 65456 526682 65512
rect 530122 57160 530178 57216
rect 529018 14456 529074 14512
rect 527822 11600 527878 11656
rect 547878 42064 547934 42120
rect 580170 72936 580226 72992
rect 577502 71848 577558 71904
rect 559746 71032 559802 71088
rect 565634 48864 565690 48920
rect 563242 29552 563298 29608
rect 564438 18672 564494 18728
rect 576122 64096 576178 64152
rect 576306 47504 576362 47560
rect 576122 6568 576178 6624
rect 577410 12960 577466 13016
rect 580722 577632 580778 577688
rect 580630 524456 580686 524512
rect 580538 208936 580594 208992
rect 580538 152632 580594 152688
rect 580446 149640 580502 149696
rect 580446 112784 580502 112840
rect 580354 71576 580410 71632
rect 580814 232328 580870 232384
rect 580722 214512 580778 214568
rect 580630 135904 580686 135960
rect 580538 71440 580594 71496
rect 580998 46144 581054 46200
rect 580262 33088 580318 33144
rect 578606 18536 578662 18592
<< metal3 >>
rect 45369 700634 45435 700637
rect 154113 700634 154179 700637
rect 45369 700632 154179 700634
rect 45369 700576 45374 700632
rect 45430 700576 154118 700632
rect 154174 700576 154179 700632
rect 45369 700574 154179 700576
rect 45369 700571 45435 700574
rect 154113 700571 154179 700574
rect 416037 700634 416103 700637
rect 429837 700634 429903 700637
rect 416037 700632 429903 700634
rect 416037 700576 416042 700632
rect 416098 700576 429842 700632
rect 429898 700576 429903 700632
rect 416037 700574 429903 700576
rect 416037 700571 416103 700574
rect 429837 700571 429903 700574
rect 44909 700498 44975 700501
rect 218973 700498 219039 700501
rect 44909 700496 219039 700498
rect 44909 700440 44914 700496
rect 44970 700440 218978 700496
rect 219034 700440 219039 700496
rect 44909 700438 219039 700440
rect 44909 700435 44975 700438
rect 218973 700435 219039 700438
rect 220077 700498 220143 700501
rect 235165 700498 235231 700501
rect 220077 700496 235231 700498
rect 220077 700440 220082 700496
rect 220138 700440 235170 700496
rect 235226 700440 235231 700496
rect 220077 700438 235231 700440
rect 220077 700435 220143 700438
rect 235165 700435 235231 700438
rect 364977 700498 365043 700501
rect 396533 700498 396599 700501
rect 364977 700496 396599 700498
rect 364977 700440 364982 700496
rect 365038 700440 396538 700496
rect 396594 700440 396599 700496
rect 364977 700438 396599 700440
rect 364977 700435 365043 700438
rect 396533 700435 396599 700438
rect 414657 700498 414723 700501
rect 494789 700498 494855 700501
rect 414657 700496 494855 700498
rect 414657 700440 414662 700496
rect 414718 700440 494794 700496
rect 494850 700440 494855 700496
rect 414657 700438 494855 700440
rect 414657 700435 414723 700438
rect 494789 700435 494855 700438
rect 45737 700362 45803 700365
rect 283833 700362 283899 700365
rect 45737 700360 283899 700362
rect 45737 700304 45742 700360
rect 45798 700304 283838 700360
rect 283894 700304 283899 700360
rect 45737 700302 283899 700304
rect 45737 700299 45803 700302
rect 283833 700299 283899 700302
rect 348785 700362 348851 700365
rect 396625 700362 396691 700365
rect 348785 700360 396691 700362
rect 348785 700304 348790 700360
rect 348846 700304 396630 700360
rect 396686 700304 396691 700360
rect 348785 700302 396691 700304
rect 348785 700299 348851 700302
rect 396625 700299 396691 700302
rect 406377 700362 406443 700365
rect 559649 700362 559715 700365
rect 406377 700360 559715 700362
rect 406377 700304 406382 700360
rect 406438 700304 559654 700360
rect 559710 700304 559715 700360
rect 406377 700302 559715 700304
rect 406377 700299 406443 700302
rect 559649 700299 559715 700302
rect 300117 699954 300183 699957
rect 303153 699954 303219 699957
rect 300117 699952 303219 699954
rect 300117 699896 300122 699952
rect 300178 699896 303158 699952
rect 303214 699896 303219 699952
rect 300117 699894 303219 699896
rect 300117 699891 300183 699894
rect 303153 699891 303219 699894
rect 303153 697506 303219 697509
rect 309777 697506 309843 697509
rect 303153 697504 309843 697506
rect -960 697220 480 697460
rect 303153 697448 303158 697504
rect 303214 697448 309782 697504
rect 309838 697448 309843 697504
rect 303153 697446 309843 697448
rect 303153 697443 303219 697446
rect 309777 697443 309843 697446
rect 580349 697234 580415 697237
rect 583520 697234 584960 697324
rect 580349 697232 584960 697234
rect 580349 697176 580354 697232
rect 580410 697176 584960 697232
rect 580349 697174 584960 697176
rect 580349 697171 580415 697174
rect 583520 697084 584960 697174
rect 309777 690162 309843 690165
rect 312537 690162 312603 690165
rect 309777 690160 312603 690162
rect 309777 690104 309782 690160
rect 309838 690104 312542 690160
rect 312598 690104 312603 690160
rect 309777 690102 312603 690104
rect 309777 690099 309843 690102
rect 312537 690099 312603 690102
rect 312537 685810 312603 685813
rect 315297 685810 315363 685813
rect 312537 685808 315363 685810
rect 312537 685752 312542 685808
rect 312598 685752 315302 685808
rect 315358 685752 315363 685808
rect 312537 685750 315363 685752
rect 312537 685747 312603 685750
rect 315297 685747 315363 685750
rect -960 684314 480 684404
rect 15837 684314 15903 684317
rect -960 684312 15903 684314
rect -960 684256 15842 684312
rect 15898 684256 15903 684312
rect -960 684254 15903 684256
rect -960 684164 480 684254
rect 15837 684251 15903 684254
rect 580533 683906 580599 683909
rect 583520 683906 584960 683996
rect 580533 683904 584960 683906
rect 580533 683848 580538 683904
rect 580594 683848 584960 683904
rect 580533 683846 584960 683848
rect 580533 683843 580599 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 26877 671258 26943 671261
rect -960 671256 26943 671258
rect -960 671200 26882 671256
rect 26938 671200 26943 671256
rect -960 671198 26943 671200
rect -960 671108 480 671198
rect 26877 671195 26943 671198
rect 544377 670714 544443 670717
rect 583520 670714 584960 670804
rect 544377 670712 584960 670714
rect 544377 670656 544382 670712
rect 544438 670656 584960 670712
rect 544377 670654 584960 670656
rect 544377 670651 544443 670654
rect 583520 670564 584960 670654
rect 315297 663914 315363 663917
rect 317413 663914 317479 663917
rect 315297 663912 317479 663914
rect 315297 663856 315302 663912
rect 315358 663856 317418 663912
rect 317474 663856 317479 663912
rect 315297 663854 317479 663856
rect 315297 663851 315363 663854
rect 317413 663851 317479 663854
rect 317413 658882 317479 658885
rect 337377 658882 337443 658885
rect 317413 658880 337443 658882
rect 317413 658824 317418 658880
rect 317474 658824 337382 658880
rect 337438 658824 337443 658880
rect 317413 658822 337443 658824
rect 317413 658819 317479 658822
rect 337377 658819 337443 658822
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect 337377 646506 337443 646509
rect 345013 646506 345079 646509
rect 337377 646504 345079 646506
rect 337377 646448 337382 646504
rect 337438 646448 345018 646504
rect 345074 646448 345079 646504
rect 337377 646446 345079 646448
rect 337377 646443 337443 646446
rect 345013 646443 345079 646446
rect -960 644996 480 645236
rect 213177 644602 213243 644605
rect 220077 644602 220143 644605
rect 213177 644600 220143 644602
rect 213177 644544 213182 644600
rect 213238 644544 220082 644600
rect 220138 644544 220143 644600
rect 213177 644542 220143 644544
rect 213177 644539 213243 644542
rect 220077 644539 220143 644542
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect 345013 639706 345079 639709
rect 348417 639706 348483 639709
rect 345013 639704 348483 639706
rect 345013 639648 345018 639704
rect 345074 639648 348422 639704
rect 348478 639648 348483 639704
rect 345013 639646 348483 639648
rect 345013 639643 345079 639646
rect 348417 639643 348483 639646
rect -960 632090 480 632180
rect 18597 632090 18663 632093
rect -960 632088 18663 632090
rect -960 632032 18602 632088
rect 18658 632032 18663 632088
rect -960 632030 18663 632032
rect -960 631940 480 632030
rect 18597 632027 18663 632030
rect 580441 630866 580507 630869
rect 583520 630866 584960 630956
rect 580441 630864 584960 630866
rect 580441 630808 580446 630864
rect 580502 630808 584960 630864
rect 580441 630806 584960 630808
rect 580441 630803 580507 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 29637 619170 29703 619173
rect -960 619168 29703 619170
rect -960 619112 29642 619168
rect 29698 619112 29703 619168
rect -960 619110 29703 619112
rect -960 619020 480 619110
rect 29637 619107 29703 619110
rect 404997 617538 405063 617541
rect 583520 617538 584960 617628
rect 404997 617536 584960 617538
rect 404997 617480 405002 617536
rect 405058 617480 584960 617536
rect 404997 617478 584960 617480
rect 404997 617475 405063 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579705 591018 579771 591021
rect 583520 591018 584960 591108
rect 579705 591016 584960 591018
rect 579705 590960 579710 591016
rect 579766 590960 584960 591016
rect 579705 590958 584960 590960
rect 579705 590955 579771 590958
rect 583520 590868 584960 590958
rect 207657 589930 207723 589933
rect 213177 589930 213243 589933
rect 207657 589928 213243 589930
rect 207657 589872 207662 589928
rect 207718 589872 213182 589928
rect 213238 589872 213243 589928
rect 207657 589870 213243 589872
rect 207657 589867 207723 589870
rect 213177 589867 213243 589870
rect -960 580002 480 580092
rect 22737 580002 22803 580005
rect -960 580000 22803 580002
rect -960 579944 22742 580000
rect 22798 579944 22803 580000
rect -960 579942 22803 579944
rect -960 579852 480 579942
rect 22737 579939 22803 579942
rect 580717 577690 580783 577693
rect 583520 577690 584960 577780
rect 580717 577688 584960 577690
rect 580717 577632 580722 577688
rect 580778 577632 584960 577688
rect 580717 577630 584960 577632
rect 580717 577627 580783 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3693 566946 3759 566949
rect -960 566944 3759 566946
rect -960 566888 3698 566944
rect 3754 566888 3759 566944
rect -960 566886 3759 566888
rect -960 566796 480 566886
rect 3693 566883 3759 566886
rect 403617 564362 403683 564365
rect 583520 564362 584960 564452
rect 403617 564360 584960 564362
rect 403617 564304 403622 564360
rect 403678 564304 584960 564360
rect 403617 564302 584960 564304
rect 403617 564299 403683 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 204897 551986 204963 551989
rect 207657 551986 207723 551989
rect 204897 551984 207723 551986
rect 204897 551928 204902 551984
rect 204958 551928 207662 551984
rect 207718 551928 207723 551984
rect 204897 551926 207723 551928
rect 204897 551923 204963 551926
rect 207657 551923 207723 551926
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 31017 527914 31083 527917
rect -960 527912 31083 527914
rect -960 527856 31022 527912
rect 31078 527856 31083 527912
rect -960 527854 31083 527856
rect -960 527764 480 527854
rect 31017 527851 31083 527854
rect 348417 525874 348483 525877
rect 351177 525874 351243 525877
rect 348417 525872 351243 525874
rect 348417 525816 348422 525872
rect 348478 525816 351182 525872
rect 351238 525816 351243 525872
rect 348417 525814 351243 525816
rect 348417 525811 348483 525814
rect 351177 525811 351243 525814
rect 580625 524514 580691 524517
rect 583520 524514 584960 524604
rect 580625 524512 584960 524514
rect 580625 524456 580630 524512
rect 580686 524456 584960 524512
rect 580625 524454 584960 524456
rect 580625 524451 580691 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 4797 514858 4863 514861
rect -960 514856 4863 514858
rect -960 514800 4802 514856
rect 4858 514800 4863 514856
rect -960 514798 4863 514800
rect -960 514708 480 514798
rect 4797 514795 4863 514798
rect 400857 511322 400923 511325
rect 583520 511322 584960 511412
rect 400857 511320 584960 511322
rect 400857 511264 400862 511320
rect 400918 511264 584960 511320
rect 400857 511262 584960 511264
rect 400857 511259 400923 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 197261 480858 197327 480861
rect 204897 480858 204963 480861
rect 197261 480856 204963 480858
rect 197261 480800 197266 480856
rect 197322 480800 204902 480856
rect 204958 480800 204963 480856
rect 197261 480798 204963 480800
rect 197261 480795 197327 480798
rect 204897 480795 204963 480798
rect 184197 478138 184263 478141
rect 197261 478138 197327 478141
rect 184197 478136 197327 478138
rect 184197 478080 184202 478136
rect 184258 478080 197266 478136
rect 197322 478080 197327 478136
rect 184197 478078 197327 478080
rect 184197 478075 184263 478078
rect 197261 478075 197327 478078
rect -960 475690 480 475780
rect 25497 475690 25563 475693
rect -960 475688 25563 475690
rect -960 475632 25502 475688
rect 25558 475632 25563 475688
rect -960 475630 25563 475632
rect -960 475540 480 475630
rect 25497 475627 25563 475630
rect 446397 471474 446463 471477
rect 583520 471474 584960 471564
rect 446397 471472 584960 471474
rect 446397 471416 446402 471472
rect 446458 471416 584960 471472
rect 446397 471414 584960 471416
rect 446397 471411 446463 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 4981 462634 5047 462637
rect -960 462632 5047 462634
rect -960 462576 4986 462632
rect 5042 462576 5047 462632
rect -960 462574 5047 462576
rect -960 462484 480 462574
rect 4981 462571 5047 462574
rect 399477 458146 399543 458149
rect 583520 458146 584960 458236
rect 399477 458144 584960 458146
rect 399477 458088 399482 458144
rect 399538 458088 584960 458144
rect 399477 458086 584960 458088
rect 399477 458083 399543 458086
rect 583520 457996 584960 458086
rect 178677 457466 178743 457469
rect 184197 457466 184263 457469
rect 178677 457464 184263 457466
rect 178677 457408 178682 457464
rect 178738 457408 184202 457464
rect 184258 457408 184263 457464
rect 178677 457406 184263 457408
rect 178677 457403 178743 457406
rect 184197 457403 184263 457406
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect 167637 440874 167703 440877
rect 178677 440874 178743 440877
rect 167637 440872 178743 440874
rect 167637 440816 167642 440872
rect 167698 440816 178682 440872
rect 178738 440816 178743 440872
rect 167637 440814 178743 440816
rect 167637 440811 167703 440814
rect 178677 440811 178743 440814
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 164877 427954 164943 427957
rect 167637 427954 167703 427957
rect 164877 427952 167703 427954
rect 164877 427896 164882 427952
rect 164938 427896 167642 427952
rect 167698 427896 167703 427952
rect 164877 427894 167703 427896
rect 164877 427891 164943 427894
rect 167637 427891 167703 427894
rect -960 423602 480 423692
rect 3601 423602 3667 423605
rect -960 423600 3667 423602
rect -960 423544 3606 423600
rect 3662 423544 3667 423600
rect -960 423542 3667 423544
rect -960 423452 480 423542
rect 3601 423539 3667 423542
rect 439497 418298 439563 418301
rect 583520 418298 584960 418388
rect 439497 418296 584960 418298
rect 439497 418240 439502 418296
rect 439558 418240 584960 418296
rect 439497 418238 584960 418240
rect 439497 418235 439563 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 11697 410546 11763 410549
rect -960 410544 11763 410546
rect -960 410488 11702 410544
rect 11758 410488 11763 410544
rect -960 410486 11763 410488
rect -960 410396 480 410486
rect 11697 410483 11763 410486
rect 411897 404970 411963 404973
rect 583520 404970 584960 405060
rect 411897 404968 584960 404970
rect 411897 404912 411902 404968
rect 411958 404912 584960 404968
rect 411897 404910 584960 404912
rect 411897 404907 411963 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 3693 384298 3759 384301
rect 25589 384298 25655 384301
rect 3693 384296 25655 384298
rect 3693 384240 3698 384296
rect 3754 384240 25594 384296
rect 25650 384240 25655 384296
rect 3693 384238 25655 384240
rect 3693 384235 3759 384238
rect 25589 384235 25655 384238
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 26969 371378 27035 371381
rect -960 371376 27035 371378
rect -960 371320 26974 371376
rect 27030 371320 27035 371376
rect -960 371318 27035 371320
rect -960 371228 480 371318
rect 26969 371315 27035 371318
rect 433977 365122 434043 365125
rect 583520 365122 584960 365212
rect 433977 365120 584960 365122
rect 433977 365064 433982 365120
rect 434038 365064 584960 365120
rect 433977 365062 584960 365064
rect 433977 365059 434043 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 14457 358458 14523 358461
rect -960 358456 14523 358458
rect -960 358400 14462 358456
rect 14518 358400 14523 358456
rect -960 358398 14523 358400
rect -960 358308 480 358398
rect 14457 358395 14523 358398
rect 153837 356690 153903 356693
rect 164877 356690 164943 356693
rect 153837 356688 164943 356690
rect 153837 356632 153842 356688
rect 153898 356632 164882 356688
rect 164938 356632 164943 356688
rect 153837 356630 164943 356632
rect 153837 356627 153903 356630
rect 164877 356627 164943 356630
rect 420177 351930 420243 351933
rect 583520 351930 584960 352020
rect 420177 351928 584960 351930
rect 420177 351872 420182 351928
rect 420238 351872 584960 351928
rect 420177 351870 584960 351872
rect 420177 351867 420243 351870
rect 583520 351780 584960 351870
rect 351177 351114 351243 351117
rect 376017 351114 376083 351117
rect 351177 351112 376083 351114
rect 351177 351056 351182 351112
rect 351238 351056 376022 351112
rect 376078 351056 376083 351112
rect 351177 351054 376083 351056
rect 351177 351051 351243 351054
rect 376017 351051 376083 351054
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 145833 342138 145899 342141
rect 153837 342138 153903 342141
rect 145833 342136 153903 342138
rect 145833 342080 145838 342136
rect 145894 342080 153842 342136
rect 153898 342080 153903 342136
rect 145833 342078 153903 342080
rect 145833 342075 145899 342078
rect 153837 342075 153903 342078
rect 376017 339418 376083 339421
rect 378777 339418 378843 339421
rect 376017 339416 378843 339418
rect 376017 339360 376022 339416
rect 376078 339360 378782 339416
rect 378838 339360 378843 339416
rect 376017 339358 378843 339360
rect 376017 339355 376083 339358
rect 378777 339355 378843 339358
rect 583520 338452 584960 338692
rect 142797 338058 142863 338061
rect 145833 338058 145899 338061
rect 142797 338056 145899 338058
rect 142797 338000 142802 338056
rect 142858 338000 145838 338056
rect 145894 338000 145899 338056
rect 142797 337998 145899 338000
rect 142797 337995 142863 337998
rect 145833 337995 145899 337998
rect 77937 334658 78003 334661
rect 170305 334658 170371 334661
rect 77937 334656 170371 334658
rect 77937 334600 77942 334656
rect 77998 334600 170310 334656
rect 170366 334600 170371 334656
rect 77937 334598 170371 334600
rect 77937 334595 78003 334598
rect 170305 334595 170371 334598
rect 378777 332482 378843 332485
rect 384573 332482 384639 332485
rect 378777 332480 384639 332482
rect -960 332196 480 332436
rect 378777 332424 378782 332480
rect 378838 332424 384578 332480
rect 384634 332424 384639 332480
rect 378777 332422 384639 332424
rect 378777 332419 378843 332422
rect 384573 332419 384639 332422
rect 384573 329082 384639 329085
rect 395337 329082 395403 329085
rect 384573 329080 395403 329082
rect 384573 329024 384578 329080
rect 384634 329024 395342 329080
rect 395398 329024 395403 329080
rect 384573 329022 395403 329024
rect 384573 329019 384639 329022
rect 395337 329019 395403 329022
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect 139393 323642 139459 323645
rect 142797 323642 142863 323645
rect 139393 323640 142863 323642
rect 139393 323584 139398 323640
rect 139454 323584 142802 323640
rect 142858 323584 142863 323640
rect 139393 323582 142863 323584
rect 139393 323579 139459 323582
rect 142797 323579 142863 323582
rect 76557 320922 76623 320925
rect 77937 320922 78003 320925
rect 76557 320920 78003 320922
rect 76557 320864 76562 320920
rect 76618 320864 77942 320920
rect 77998 320864 78003 320920
rect 76557 320862 78003 320864
rect 76557 320859 76623 320862
rect 77937 320859 78003 320862
rect -960 319290 480 319380
rect 29729 319290 29795 319293
rect -960 319288 29795 319290
rect -960 319232 29734 319288
rect 29790 319232 29795 319288
rect -960 319230 29795 319232
rect -960 319140 480 319230
rect 29729 319227 29795 319230
rect 128997 316706 129063 316709
rect 139393 316706 139459 316709
rect 128997 316704 139459 316706
rect 128997 316648 129002 316704
rect 129058 316648 139398 316704
rect 139454 316648 139459 316704
rect 128997 316646 139459 316648
rect 128997 316643 129063 316646
rect 139393 316643 139459 316646
rect 438117 312082 438183 312085
rect 583520 312082 584960 312172
rect 438117 312080 584960 312082
rect 438117 312024 438122 312080
rect 438178 312024 584960 312080
rect 438117 312022 584960 312024
rect 438117 312019 438183 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 31109 306234 31175 306237
rect -960 306232 31175 306234
rect -960 306176 31114 306232
rect 31170 306176 31175 306232
rect -960 306174 31175 306176
rect -960 306084 480 306174
rect 31109 306171 31175 306174
rect 126237 301610 126303 301613
rect 128997 301610 129063 301613
rect 126237 301608 129063 301610
rect 126237 301552 126242 301608
rect 126298 301552 129002 301608
rect 129058 301552 129063 301608
rect 126237 301550 129063 301552
rect 126237 301547 126303 301550
rect 128997 301547 129063 301550
rect 409137 298754 409203 298757
rect 583520 298754 584960 298844
rect 409137 298752 584960 298754
rect 409137 298696 409142 298752
rect 409198 298696 584960 298752
rect 409137 298694 584960 298696
rect 409137 298691 409203 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 75269 291138 75335 291141
rect 76557 291138 76623 291141
rect 75269 291136 76623 291138
rect 75269 291080 75274 291136
rect 75330 291080 76562 291136
rect 76618 291080 76623 291136
rect 75269 291078 76623 291080
rect 75269 291075 75335 291078
rect 76557 291075 76623 291078
rect 73245 288554 73311 288557
rect 75269 288554 75335 288557
rect 73245 288552 75335 288554
rect 73245 288496 73250 288552
rect 73306 288496 75274 288552
rect 75330 288496 75335 288552
rect 73245 288494 75335 288496
rect 73245 288491 73311 288494
rect 75269 288491 75335 288494
rect 120809 287738 120875 287741
rect 126237 287738 126303 287741
rect 120809 287736 126303 287738
rect 120809 287680 120814 287736
rect 120870 287680 126242 287736
rect 126298 287680 126303 287736
rect 120809 287678 126303 287680
rect 120809 287675 120875 287678
rect 126237 287675 126303 287678
rect 395337 285698 395403 285701
rect 396441 285698 396507 285701
rect 395337 285696 396507 285698
rect 395337 285640 395342 285696
rect 395398 285640 396446 285696
rect 396502 285640 396507 285696
rect 395337 285638 396507 285640
rect 395337 285635 395403 285638
rect 396441 285635 396507 285638
rect 583520 285276 584960 285516
rect 117957 282298 118023 282301
rect 120809 282298 120875 282301
rect 117957 282296 120875 282298
rect 117957 282240 117962 282296
rect 118018 282240 120814 282296
rect 120870 282240 120875 282296
rect 117957 282238 120875 282240
rect 117957 282235 118023 282238
rect 120809 282235 120875 282238
rect 70945 281618 71011 281621
rect 73245 281618 73311 281621
rect 70945 281616 73311 281618
rect 70945 281560 70950 281616
rect 71006 281560 73250 281616
rect 73306 281560 73311 281616
rect 70945 281558 73311 281560
rect 70945 281555 71011 281558
rect 73245 281555 73311 281558
rect -960 279972 480 280212
rect 69657 280122 69723 280125
rect 70945 280122 71011 280125
rect 69657 280120 71011 280122
rect 69657 280064 69662 280120
rect 69718 280064 70950 280120
rect 71006 280064 71011 280120
rect 69657 280062 71011 280064
rect 69657 280059 69723 280062
rect 70945 280059 71011 280062
rect 67817 276042 67883 276045
rect 69657 276042 69723 276045
rect 67817 276040 69723 276042
rect 67817 275984 67822 276040
rect 67878 275984 69662 276040
rect 69718 275984 69723 276040
rect 67817 275982 69723 275984
rect 67817 275979 67883 275982
rect 69657 275979 69723 275982
rect 113817 272234 113883 272237
rect 117957 272234 118023 272237
rect 113817 272232 118023 272234
rect 113817 272176 113822 272232
rect 113878 272176 117962 272232
rect 118018 272176 118023 272232
rect 113817 272174 118023 272176
rect 113817 272171 113883 272174
rect 117957 272171 118023 272174
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect 66529 270466 66595 270469
rect 67817 270466 67883 270469
rect 66529 270464 67883 270466
rect 66529 270408 66534 270464
rect 66590 270408 67822 270464
rect 67878 270408 67883 270464
rect 66529 270406 67883 270408
rect 66529 270403 66595 270406
rect 67817 270403 67883 270406
rect -960 267202 480 267292
rect 3693 267202 3759 267205
rect -960 267200 3759 267202
rect -960 267144 3698 267200
rect 3754 267144 3759 267200
rect -960 267142 3759 267144
rect -960 267052 480 267142
rect 3693 267139 3759 267142
rect 108297 266386 108363 266389
rect 113817 266386 113883 266389
rect 108297 266384 113883 266386
rect 108297 266328 108302 266384
rect 108358 266328 113822 266384
rect 113878 266328 113883 266384
rect 108297 266326 113883 266328
rect 108297 266323 108363 266326
rect 113817 266323 113883 266326
rect 65517 265026 65583 265029
rect 66529 265026 66595 265029
rect 65517 265024 66595 265026
rect 65517 264968 65522 265024
rect 65578 264968 66534 265024
rect 66590 264968 66595 265024
rect 65517 264966 66595 264968
rect 65517 264963 65583 264966
rect 66529 264963 66595 264966
rect 429837 258906 429903 258909
rect 583520 258906 584960 258996
rect 429837 258904 584960 258906
rect 429837 258848 429842 258904
rect 429898 258848 584960 258904
rect 429837 258846 584960 258848
rect 429837 258843 429903 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 22829 254146 22895 254149
rect -960 254144 22895 254146
rect -960 254088 22834 254144
rect 22890 254088 22895 254144
rect -960 254086 22895 254088
rect -960 253996 480 254086
rect 22829 254083 22895 254086
rect 105537 254010 105603 254013
rect 108297 254010 108363 254013
rect 105537 254008 108363 254010
rect 105537 253952 105542 254008
rect 105598 253952 108302 254008
rect 108358 253952 108363 254008
rect 105537 253950 108363 253952
rect 105537 253947 105603 253950
rect 108297 253947 108363 253950
rect 64137 248434 64203 248437
rect 65517 248434 65583 248437
rect 64137 248432 65583 248434
rect 64137 248376 64142 248432
rect 64198 248376 65522 248432
rect 65578 248376 65583 248432
rect 64137 248374 65583 248376
rect 64137 248371 64203 248374
rect 65517 248371 65583 248374
rect 407757 245578 407823 245581
rect 583520 245578 584960 245668
rect 407757 245576 584960 245578
rect 407757 245520 407762 245576
rect 407818 245520 584960 245576
rect 407757 245518 584960 245520
rect 407757 245515 407823 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 98913 236738 98979 236741
rect 105537 236738 105603 236741
rect 98913 236736 105603 236738
rect 98913 236680 98918 236736
rect 98974 236680 105542 236736
rect 105598 236680 105603 236736
rect 98913 236678 105603 236680
rect 98913 236675 98979 236678
rect 105537 236675 105603 236678
rect 580809 232386 580875 232389
rect 583520 232386 584960 232476
rect 580809 232384 584960 232386
rect 580809 232328 580814 232384
rect 580870 232328 584960 232384
rect 580809 232326 584960 232328
rect 580809 232323 580875 232326
rect 583520 232236 584960 232326
rect 53833 231162 53899 231165
rect 64137 231162 64203 231165
rect 53833 231160 64203 231162
rect 53833 231104 53838 231160
rect 53894 231104 64142 231160
rect 64198 231104 64203 231160
rect 53833 231102 64203 231104
rect 53833 231099 53899 231102
rect 64137 231099 64203 231102
rect 95233 230482 95299 230485
rect 98913 230482 98979 230485
rect 95233 230480 98979 230482
rect 95233 230424 95238 230480
rect 95294 230424 98918 230480
rect 98974 230424 98979 230480
rect 95233 230422 98979 230424
rect 95233 230419 95299 230422
rect 98913 230419 98979 230422
rect -960 227884 480 228124
rect 68921 226266 68987 226269
rect 105445 226266 105511 226269
rect 64830 226206 68754 226266
rect 45093 226130 45159 226133
rect 64830 226130 64890 226206
rect 45093 226128 64890 226130
rect 45093 226072 45098 226128
rect 45154 226072 64890 226128
rect 45093 226070 64890 226072
rect 68694 226130 68754 226206
rect 68921 226264 105511 226266
rect 68921 226208 68926 226264
rect 68982 226208 105450 226264
rect 105506 226208 105511 226264
rect 68921 226206 105511 226208
rect 68921 226203 68987 226206
rect 105445 226203 105511 226206
rect 89161 226130 89227 226133
rect 68694 226128 89227 226130
rect 68694 226072 89166 226128
rect 89222 226072 89227 226128
rect 68694 226070 89227 226072
rect 45093 226067 45159 226070
rect 89161 226067 89227 226070
rect 53833 225042 53899 225045
rect 48270 225040 53899 225042
rect 48270 224984 53838 225040
rect 53894 224984 53899 225040
rect 48270 224982 53899 224984
rect 45829 224906 45895 224909
rect 48270 224906 48330 224982
rect 53833 224979 53899 224982
rect 45829 224904 48330 224906
rect 45829 224848 45834 224904
rect 45890 224848 48330 224904
rect 45829 224846 48330 224848
rect 45829 224843 45895 224846
rect 44725 224226 44791 224229
rect 95233 224226 95299 224229
rect 44725 224224 95299 224226
rect 44725 224168 44730 224224
rect 44786 224168 95238 224224
rect 95294 224168 95299 224224
rect 44725 224166 95299 224168
rect 44725 224163 44791 224166
rect 95233 224163 95299 224166
rect 399569 219058 399635 219061
rect 583520 219058 584960 219148
rect 399569 219056 584960 219058
rect 399569 219000 399574 219056
rect 399630 219000 584960 219056
rect 399569 218998 584960 219000
rect 399569 218995 399635 218998
rect 583520 218908 584960 218998
rect 44725 216202 44791 216205
rect 46841 216202 46907 216205
rect 44725 216200 46907 216202
rect 44725 216144 44730 216200
rect 44786 216144 46846 216200
rect 46902 216144 46907 216200
rect 44725 216142 46907 216144
rect 44725 216139 44791 216142
rect 46841 216139 46907 216142
rect 45829 215930 45895 215933
rect 149053 215930 149119 215933
rect 45829 215928 149119 215930
rect 45829 215872 45834 215928
rect 45890 215872 149058 215928
rect 149114 215872 149119 215928
rect 45829 215870 149119 215872
rect 45829 215867 45895 215870
rect 149053 215867 149119 215870
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 3601 214842 3667 214845
rect 177849 214842 177915 214845
rect 3601 214840 177915 214842
rect 3601 214784 3606 214840
rect 3662 214784 177854 214840
rect 177910 214784 177915 214840
rect 3601 214782 177915 214784
rect 3601 214779 3667 214782
rect 177849 214779 177915 214782
rect 390553 214842 390619 214845
rect 396441 214842 396507 214845
rect 390553 214840 396507 214842
rect 390553 214784 390558 214840
rect 390614 214784 396446 214840
rect 396502 214784 396507 214840
rect 390553 214782 396507 214784
rect 390553 214779 390619 214782
rect 396441 214779 396507 214782
rect 114369 214706 114435 214709
rect 396625 214706 396691 214709
rect 114369 214704 396691 214706
rect 114369 214648 114374 214704
rect 114430 214648 396630 214704
rect 396686 214648 396691 214704
rect 114369 214646 396691 214648
rect 114369 214643 114435 214646
rect 396625 214643 396691 214646
rect 115841 214570 115907 214573
rect 580717 214570 580783 214573
rect 115841 214568 580783 214570
rect 115841 214512 115846 214568
rect 115902 214512 580722 214568
rect 580778 214512 580783 214568
rect 115841 214510 580783 214512
rect 115841 214507 115907 214510
rect 580717 214507 580783 214510
rect 149053 213210 149119 213213
rect 159357 213210 159423 213213
rect 149053 213208 159423 213210
rect 149053 213152 149058 213208
rect 149114 213152 159362 213208
rect 159418 213152 159423 213208
rect 149053 213150 159423 213152
rect 149053 213147 149119 213150
rect 159357 213147 159423 213150
rect 162117 213210 162183 213213
rect 296713 213210 296779 213213
rect 162117 213208 296779 213210
rect 162117 213152 162122 213208
rect 162178 213152 296718 213208
rect 296774 213152 296779 213208
rect 162117 213150 296779 213152
rect 162117 213147 162183 213150
rect 296713 213147 296779 213150
rect 358077 213210 358143 213213
rect 386505 213210 386571 213213
rect 358077 213208 386571 213210
rect 358077 213152 358082 213208
rect 358138 213152 386510 213208
rect 386566 213152 386571 213208
rect 358077 213150 386571 213152
rect 358077 213147 358143 213150
rect 386505 213147 386571 213150
rect 355317 212666 355383 212669
rect 356513 212666 356579 212669
rect 355317 212664 356579 212666
rect 355317 212608 355322 212664
rect 355378 212608 356518 212664
rect 356574 212608 356579 212664
rect 355317 212606 356579 212608
rect 355317 212603 355383 212606
rect 356513 212603 356579 212606
rect 3693 211850 3759 211853
rect 176837 211850 176903 211853
rect 3693 211848 176903 211850
rect 3693 211792 3698 211848
rect 3754 211792 176842 211848
rect 176898 211792 176903 211848
rect 3693 211790 176903 211792
rect 3693 211787 3759 211790
rect 176837 211787 176903 211790
rect 387333 211170 387399 211173
rect 390461 211170 390527 211173
rect 387333 211168 390527 211170
rect 387333 211112 387338 211168
rect 387394 211112 390466 211168
rect 390522 211112 390527 211168
rect 387333 211110 390527 211112
rect 387333 211107 387399 211110
rect 390461 211107 390527 211110
rect 46841 210490 46907 210493
rect 56593 210490 56659 210493
rect 46841 210488 56659 210490
rect 46841 210432 46846 210488
rect 46902 210432 56598 210488
rect 56654 210432 56659 210488
rect 46841 210430 56659 210432
rect 46841 210427 46907 210430
rect 56593 210427 56659 210430
rect 3325 210354 3391 210357
rect 175273 210354 175339 210357
rect 3325 210352 175339 210354
rect 3325 210296 3330 210352
rect 3386 210296 175278 210352
rect 175334 210296 175339 210352
rect 3325 210294 175339 210296
rect 3325 210291 3391 210294
rect 175273 210291 175339 210294
rect 159357 209130 159423 209133
rect 167637 209130 167703 209133
rect 159357 209128 167703 209130
rect 159357 209072 159362 209128
rect 159418 209072 167642 209128
rect 167698 209072 167703 209128
rect 159357 209070 167703 209072
rect 159357 209067 159423 209070
rect 167637 209067 167703 209070
rect 115749 208994 115815 208997
rect 580533 208994 580599 208997
rect 115749 208992 580599 208994
rect 115749 208936 115754 208992
rect 115810 208936 580538 208992
rect 580594 208936 580599 208992
rect 115749 208934 580599 208936
rect 115749 208931 115815 208934
rect 580533 208931 580599 208934
rect 383653 208450 383719 208453
rect 387333 208450 387399 208453
rect 383653 208448 387399 208450
rect 383653 208392 383658 208448
rect 383714 208392 387338 208448
rect 387394 208392 387399 208448
rect 383653 208390 387399 208392
rect 383653 208387 383719 208390
rect 387333 208387 387399 208390
rect 143441 207090 143507 207093
rect 146293 207090 146359 207093
rect 143441 207088 146359 207090
rect 143441 207032 143446 207088
rect 143502 207032 146298 207088
rect 146354 207032 146359 207088
rect 143441 207030 146359 207032
rect 143441 207027 143507 207030
rect 146293 207027 146359 207030
rect 56593 205730 56659 205733
rect 58617 205730 58683 205733
rect 56593 205728 58683 205730
rect 56593 205672 56598 205728
rect 56654 205672 58622 205728
rect 58678 205672 58683 205728
rect 56593 205670 58683 205672
rect 56593 205667 56659 205670
rect 58617 205667 58683 205670
rect 188337 205730 188403 205733
rect 583520 205730 584960 205820
rect 188337 205728 584960 205730
rect 188337 205672 188342 205728
rect 188398 205672 584960 205728
rect 188337 205670 584960 205672
rect 188337 205667 188403 205670
rect 583520 205580 584960 205670
rect 378133 204370 378199 204373
rect 383561 204370 383627 204373
rect 378133 204368 383627 204370
rect 378133 204312 378138 204368
rect 378194 204312 383566 204368
rect 383622 204312 383627 204368
rect 378133 204310 383627 204312
rect 378133 204307 378199 204310
rect 383561 204307 383627 204310
rect 114461 203554 114527 203557
rect 399569 203554 399635 203557
rect 114461 203552 399635 203554
rect 114461 203496 114466 203552
rect 114522 203496 399574 203552
rect 399630 203496 399635 203552
rect 114461 203494 399635 203496
rect 114461 203491 114527 203494
rect 399569 203491 399635 203494
rect -960 201922 480 202012
rect 46197 201922 46263 201925
rect -960 201920 46263 201922
rect -960 201864 46202 201920
rect 46258 201864 46263 201920
rect -960 201862 46263 201864
rect -960 201772 480 201862
rect 46197 201859 46263 201862
rect 375373 201378 375439 201381
rect 378041 201378 378107 201381
rect 375373 201376 378107 201378
rect 375373 201320 375378 201376
rect 375434 201320 378046 201376
rect 378102 201320 378107 201376
rect 375373 201318 378107 201320
rect 375373 201315 375439 201318
rect 378041 201315 378107 201318
rect 167637 198794 167703 198797
rect 173157 198794 173223 198797
rect 375373 198794 375439 198797
rect 167637 198792 173223 198794
rect 167637 198736 167642 198792
rect 167698 198736 173162 198792
rect 173218 198736 173223 198792
rect 167637 198734 173223 198736
rect 167637 198731 167703 198734
rect 173157 198731 173223 198734
rect 373950 198792 375439 198794
rect 373950 198736 375378 198792
rect 375434 198736 375439 198792
rect 373950 198734 375439 198736
rect 369853 198658 369919 198661
rect 373950 198658 374010 198734
rect 375373 198731 375439 198734
rect 369853 198656 374010 198658
rect 369853 198600 369858 198656
rect 369914 198600 374010 198656
rect 369853 198598 374010 198600
rect 369853 198595 369919 198598
rect 116761 195258 116827 195261
rect 478505 195258 478571 195261
rect 116761 195256 478571 195258
rect 116761 195200 116766 195256
rect 116822 195200 478510 195256
rect 478566 195200 478571 195256
rect 116761 195198 478571 195200
rect 116761 195195 116827 195198
rect 478505 195195 478571 195198
rect 57881 193898 57947 193901
rect 134517 193898 134583 193901
rect 57881 193896 134583 193898
rect 57881 193840 57886 193896
rect 57942 193840 134522 193896
rect 134578 193840 134583 193896
rect 57881 193838 134583 193840
rect 57881 193835 57947 193838
rect 134517 193835 134583 193838
rect 363597 193898 363663 193901
rect 369761 193898 369827 193901
rect 363597 193896 369827 193898
rect 363597 193840 363602 193896
rect 363658 193840 369766 193896
rect 369822 193840 369827 193896
rect 363597 193838 369827 193840
rect 363597 193835 363663 193838
rect 369761 193835 369827 193838
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 58617 191722 58683 191725
rect 59997 191722 60063 191725
rect 58617 191720 60063 191722
rect 58617 191664 58622 191720
rect 58678 191664 60002 191720
rect 60058 191664 60063 191720
rect 58617 191662 60063 191664
rect 58617 191659 58683 191662
rect 59997 191659 60063 191662
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 157241 186962 157307 186965
rect 355317 186962 355383 186965
rect 157241 186960 355383 186962
rect 157241 186904 157246 186960
rect 157302 186904 355322 186960
rect 355378 186904 355383 186960
rect 157241 186902 355383 186904
rect 157241 186899 157307 186902
rect 355317 186899 355383 186902
rect 59997 186418 60063 186421
rect 61377 186418 61443 186421
rect 59997 186416 61443 186418
rect 59997 186360 60002 186416
rect 60058 186360 61382 186416
rect 61438 186360 61443 186416
rect 59997 186358 61443 186360
rect 59997 186355 60063 186358
rect 61377 186355 61443 186358
rect 173157 186418 173223 186421
rect 175917 186418 175983 186421
rect 173157 186416 175983 186418
rect 173157 186360 173162 186416
rect 173218 186360 175922 186416
rect 175978 186360 175983 186416
rect 173157 186358 175983 186360
rect 173157 186355 173223 186358
rect 175917 186355 175983 186358
rect 360837 186418 360903 186421
rect 363597 186418 363663 186421
rect 360837 186416 363663 186418
rect 360837 186360 360842 186416
rect 360898 186360 363602 186416
rect 363658 186360 363663 186416
rect 360837 186358 363663 186360
rect 360837 186355 360903 186358
rect 363597 186355 363663 186358
rect 152733 184242 152799 184245
rect 327073 184242 327139 184245
rect 152733 184240 327139 184242
rect 152733 184184 152738 184240
rect 152794 184184 327078 184240
rect 327134 184184 327139 184240
rect 152733 184182 327139 184184
rect 152733 184179 152799 184182
rect 327073 184179 327139 184182
rect 155953 183562 156019 183565
rect 358077 183562 358143 183565
rect 155953 183560 358143 183562
rect 155953 183504 155958 183560
rect 156014 183504 358082 183560
rect 358138 183504 358143 183560
rect 155953 183502 358143 183504
rect 155953 183499 156019 183502
rect 358077 183499 358143 183502
rect 154297 183426 154363 183429
rect 157241 183426 157307 183429
rect 154297 183424 157307 183426
rect 154297 183368 154302 183424
rect 154358 183368 157246 183424
rect 157302 183368 157307 183424
rect 154297 183366 157307 183368
rect 154297 183363 154363 183366
rect 157241 183363 157307 183366
rect 88241 182066 88307 182069
rect 133229 182066 133295 182069
rect 88241 182064 133295 182066
rect 88241 182008 88246 182064
rect 88302 182008 133234 182064
rect 133290 182008 133295 182064
rect 88241 182006 133295 182008
rect 88241 182003 88307 182006
rect 133229 182003 133295 182006
rect 136633 182066 136699 182069
rect 136633 182064 139042 182066
rect 136633 182008 136638 182064
rect 136694 182008 139042 182064
rect 136633 182006 139042 182008
rect 136633 182003 136699 182006
rect 138982 181998 139042 182006
rect 138982 181938 139564 181998
rect 155769 181794 155835 181797
rect 162117 181794 162183 181797
rect 155769 181792 162183 181794
rect 155769 181736 155774 181792
rect 155830 181736 162122 181792
rect 162178 181736 162183 181792
rect 155769 181734 162183 181736
rect 155769 181731 155835 181734
rect 162117 181731 162183 181734
rect 138565 181386 138631 181389
rect 137970 181384 138631 181386
rect 137970 181328 138570 181384
rect 138626 181328 138631 181384
rect 137970 181326 138631 181328
rect 137829 181250 137895 181253
rect 137970 181250 138030 181326
rect 138565 181323 138631 181326
rect 154481 181386 154547 181389
rect 155401 181386 155467 181389
rect 154481 181384 155467 181386
rect 154481 181328 154486 181384
rect 154542 181328 155406 181384
rect 155462 181328 155467 181384
rect 154481 181326 155467 181328
rect 154481 181323 154547 181326
rect 155401 181323 155467 181326
rect 163037 181386 163103 181389
rect 442257 181386 442323 181389
rect 163037 181384 442323 181386
rect 163037 181328 163042 181384
rect 163098 181328 442262 181384
rect 442318 181328 442323 181384
rect 163037 181326 442323 181328
rect 163037 181323 163103 181326
rect 442257 181323 442323 181326
rect 138749 181250 138815 181253
rect 137829 181248 138030 181250
rect 137829 181192 137834 181248
rect 137890 181192 138030 181248
rect 137829 181190 138030 181192
rect 138246 181248 138815 181250
rect 138246 181192 138754 181248
rect 138810 181192 138815 181248
rect 138246 181190 138815 181192
rect 137829 181187 137895 181190
rect 136030 181052 136036 181116
rect 136100 181114 136106 181116
rect 138013 181114 138079 181117
rect 136100 181112 138079 181114
rect 136100 181056 138018 181112
rect 138074 181056 138079 181112
rect 136100 181054 138079 181056
rect 136100 181052 136106 181054
rect 138013 181051 138079 181054
rect 135846 180916 135852 180980
rect 135916 180978 135922 180980
rect 138246 180978 138306 181190
rect 138749 181187 138815 181190
rect 135916 180918 138306 180978
rect 135916 180916 135922 180918
rect 117221 180706 117287 180709
rect 133229 180706 133295 180709
rect 117221 180704 133295 180706
rect 117221 180648 117226 180704
rect 117282 180648 133234 180704
rect 133290 180648 133295 180704
rect 117221 180646 133295 180648
rect 117221 180643 117287 180646
rect 133229 180643 133295 180646
rect 140957 179754 141023 179757
rect 143950 179754 144010 180264
rect 149881 180026 149947 180029
rect 155401 180026 155467 180029
rect 149881 180024 155467 180026
rect 149881 179968 149886 180024
rect 149942 179968 155406 180024
rect 155462 179968 155467 180024
rect 149881 179966 155467 179968
rect 149881 179963 149947 179966
rect 155401 179963 155467 179966
rect 151721 179890 151787 179893
rect 155493 179890 155559 179893
rect 151721 179888 155559 179890
rect 151721 179832 151726 179888
rect 151782 179832 155498 179888
rect 155554 179832 155559 179888
rect 151721 179830 155559 179832
rect 151721 179827 151787 179830
rect 155493 179827 155559 179830
rect 140957 179752 144010 179754
rect 140957 179696 140962 179752
rect 141018 179696 144010 179752
rect 140957 179694 144010 179696
rect 150985 179754 151051 179757
rect 155769 179754 155835 179757
rect 150985 179752 155835 179754
rect 150985 179696 150990 179752
rect 151046 179696 155774 179752
rect 155830 179696 155835 179752
rect 150985 179694 155835 179696
rect 140957 179691 141023 179694
rect 150985 179691 151051 179694
rect 155769 179691 155835 179694
rect 146017 179618 146083 179621
rect 137970 179616 146083 179618
rect 137970 179560 146022 179616
rect 146078 179560 146083 179616
rect 137970 179558 146083 179560
rect 136357 179482 136423 179485
rect 137970 179482 138030 179558
rect 146017 179555 146083 179558
rect 136357 179480 138030 179482
rect 136357 179424 136362 179480
rect 136418 179424 138030 179480
rect 136357 179422 138030 179424
rect 146293 179482 146359 179485
rect 162761 179482 162827 179485
rect 146293 179480 162827 179482
rect 146293 179424 146298 179480
rect 146354 179424 162766 179480
rect 162822 179424 162827 179480
rect 146293 179422 162827 179424
rect 136357 179419 136423 179422
rect 146293 179419 146359 179422
rect 162761 179419 162827 179422
rect 199377 179210 199443 179213
rect 583520 179210 584960 179300
rect 199377 179208 584960 179210
rect 199377 179152 199382 179208
rect 199438 179152 584960 179208
rect 199377 179150 584960 179152
rect 199377 179147 199443 179150
rect 583520 179060 584960 179150
rect 140630 178068 140636 178132
rect 140700 178130 140706 178132
rect 140700 178070 141220 178130
rect 140700 178068 140706 178070
rect 139526 177380 139532 177444
rect 139596 177442 139602 177444
rect 141190 177442 141250 177960
rect 139596 177382 141250 177442
rect 139596 177380 139602 177382
rect -960 175796 480 176036
rect 141918 176020 141924 176084
rect 141988 176082 141994 176084
rect 142613 176082 142679 176085
rect 141988 176080 142679 176082
rect 141988 176024 142618 176080
rect 142674 176024 142679 176080
rect 141988 176022 142679 176024
rect 141988 176020 141994 176022
rect 142613 176019 142679 176022
rect 359457 173906 359523 173909
rect 360837 173906 360903 173909
rect 359457 173904 360903 173906
rect 359457 173848 359462 173904
rect 359518 173848 360842 173904
rect 360898 173848 360903 173904
rect 359457 173846 360903 173848
rect 359457 173843 359523 173846
rect 360837 173843 360903 173846
rect 141550 172484 141556 172548
rect 141620 172546 141626 172548
rect 141877 172546 141943 172549
rect 141620 172544 141943 172546
rect 141620 172488 141882 172544
rect 141938 172488 141943 172544
rect 141620 172486 141943 172488
rect 141620 172484 141626 172486
rect 141877 172483 141943 172486
rect 61377 167106 61443 167109
rect 62757 167106 62823 167109
rect 61377 167104 62823 167106
rect 61377 167048 61382 167104
rect 61438 167048 62762 167104
rect 62818 167048 62823 167104
rect 61377 167046 62823 167048
rect 61377 167043 61443 167046
rect 62757 167043 62823 167046
rect 185577 165882 185643 165885
rect 583520 165882 584960 165972
rect 185577 165880 584960 165882
rect 185577 165824 185582 165880
rect 185638 165824 584960 165880
rect 185577 165822 584960 165824
rect 185577 165819 185643 165822
rect 583520 165732 584960 165822
rect 139485 165204 139551 165205
rect 139485 165202 139532 165204
rect 139440 165200 139532 165202
rect 139440 165144 139490 165200
rect 139440 165142 139532 165144
rect 139485 165140 139532 165142
rect 139596 165140 139602 165204
rect 139485 165139 139551 165140
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 141550 162148 141556 162212
rect 141620 162210 141626 162212
rect 168373 162210 168439 162213
rect 141620 162208 168439 162210
rect 141620 162152 168378 162208
rect 168434 162152 168439 162208
rect 141620 162150 168439 162152
rect 141620 162148 141626 162150
rect 168373 162147 168439 162150
rect 3325 162074 3391 162077
rect 136081 162074 136147 162077
rect 3325 162072 136147 162074
rect 3325 162016 3330 162072
rect 3386 162016 136086 162072
rect 136142 162016 136147 162072
rect 3325 162014 136147 162016
rect 3325 162011 3391 162014
rect 136081 162011 136147 162014
rect 136357 162074 136423 162077
rect 176745 162074 176811 162077
rect 136357 162072 176811 162074
rect 136357 162016 136362 162072
rect 136418 162016 176750 162072
rect 176806 162016 176811 162072
rect 136357 162014 176811 162016
rect 136357 162011 136423 162014
rect 176745 162011 176811 162014
rect 135846 161530 135852 161532
rect 135302 161470 135852 161530
rect 135302 160034 135362 161470
rect 135846 161468 135852 161470
rect 135916 161468 135922 161532
rect 160461 161530 160527 161533
rect 163221 161530 163287 161533
rect 160461 161528 163287 161530
rect 160461 161472 160466 161528
rect 160522 161472 163226 161528
rect 163282 161472 163287 161528
rect 160461 161470 163287 161472
rect 160461 161467 160527 161470
rect 163221 161467 163287 161470
rect 136398 161332 136404 161396
rect 136468 161332 136474 161396
rect 135846 160034 135852 160036
rect 135302 159974 135852 160034
rect 135846 159972 135852 159974
rect 135916 159972 135922 160036
rect 136030 159972 136036 160036
rect 136100 160034 136106 160036
rect 136406 160034 136466 161332
rect 139485 161122 139551 161125
rect 139485 161120 142170 161122
rect 139485 161064 139490 161120
rect 139546 161064 142170 161120
rect 139485 161062 142170 161064
rect 139485 161059 139551 161062
rect 142110 160714 142170 161062
rect 163681 160714 163747 160717
rect 142110 160712 163747 160714
rect 142110 160656 163686 160712
rect 163742 160656 163747 160712
rect 142110 160654 163747 160656
rect 163681 160651 163747 160654
rect 136100 159974 136466 160034
rect 136100 159972 136106 159974
rect 114001 156634 114067 156637
rect 433977 156634 434043 156637
rect 114001 156632 434043 156634
rect 114001 156576 114006 156632
rect 114062 156576 433982 156632
rect 434038 156576 434043 156632
rect 114001 156574 434043 156576
rect 114001 156571 114067 156574
rect 433977 156571 434043 156574
rect 114093 155274 114159 155277
rect 438117 155274 438183 155277
rect 114093 155272 438183 155274
rect 114093 155216 114098 155272
rect 114154 155216 438122 155272
rect 438178 155216 438183 155272
rect 114093 155214 438183 155216
rect 114093 155211 114159 155214
rect 438117 155211 438183 155214
rect 114185 153778 114251 153781
rect 429837 153778 429903 153781
rect 114185 153776 429903 153778
rect 114185 153720 114190 153776
rect 114246 153720 429842 153776
rect 429898 153720 429903 153776
rect 114185 153718 429903 153720
rect 114185 153715 114251 153718
rect 429837 153715 429903 153718
rect 580533 152690 580599 152693
rect 583520 152690 584960 152780
rect 580533 152688 584960 152690
rect 580533 152632 580538 152688
rect 580594 152632 584960 152688
rect 580533 152630 584960 152632
rect 580533 152627 580599 152630
rect 583520 152540 584960 152630
rect 140630 152356 140636 152420
rect 140700 152418 140706 152420
rect 161565 152418 161631 152421
rect 140700 152416 161631 152418
rect 140700 152360 161570 152416
rect 161626 152360 161631 152416
rect 140700 152358 161631 152360
rect 140700 152356 140706 152358
rect 161565 152355 161631 152358
rect 114277 151058 114343 151061
rect 199377 151058 199443 151061
rect 114277 151056 199443 151058
rect 114277 151000 114282 151056
rect 114338 151000 199382 151056
rect 199438 151000 199443 151056
rect 114277 150998 199443 151000
rect 114277 150995 114343 150998
rect 199377 150995 199443 150998
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 115657 149698 115723 149701
rect 580441 149698 580507 149701
rect 115657 149696 580507 149698
rect 115657 149640 115662 149696
rect 115718 149640 580446 149696
rect 580502 149640 580507 149696
rect 115657 149638 580507 149640
rect 115657 149635 115723 149638
rect 580441 149635 580507 149638
rect 355685 149154 355751 149157
rect 359457 149154 359523 149157
rect 355685 149152 359523 149154
rect 355685 149096 355690 149152
rect 355746 149096 359462 149152
rect 359518 149096 359523 149152
rect 355685 149094 359523 149096
rect 355685 149091 355751 149094
rect 359457 149091 359523 149094
rect 29729 148338 29795 148341
rect 178769 148338 178835 148341
rect 29729 148336 178835 148338
rect 29729 148280 29734 148336
rect 29790 148280 178774 148336
rect 178830 148280 178835 148336
rect 29729 148278 178835 148280
rect 29729 148275 29795 148278
rect 178769 148275 178835 148278
rect 26969 146978 27035 146981
rect 178677 146978 178743 146981
rect 26969 146976 178743 146978
rect 26969 146920 26974 146976
rect 27030 146920 178682 146976
rect 178738 146920 178743 146976
rect 26969 146918 178743 146920
rect 26969 146915 27035 146918
rect 178677 146915 178743 146918
rect 25497 145618 25563 145621
rect 178217 145618 178283 145621
rect 25497 145616 178283 145618
rect 25497 145560 25502 145616
rect 25558 145560 178222 145616
rect 178278 145560 178283 145616
rect 25497 145558 178283 145560
rect 25497 145555 25563 145558
rect 178217 145555 178283 145558
rect 62757 144258 62823 144261
rect 70761 144258 70827 144261
rect 62757 144256 70827 144258
rect 62757 144200 62762 144256
rect 62818 144200 70766 144256
rect 70822 144200 70827 144256
rect 62757 144198 70827 144200
rect 62757 144195 62823 144198
rect 70761 144195 70827 144198
rect 31017 144122 31083 144125
rect 178309 144122 178375 144125
rect 31017 144120 178375 144122
rect 31017 144064 31022 144120
rect 31078 144064 178314 144120
rect 178370 144064 178375 144120
rect 31017 144062 178375 144064
rect 31017 144059 31083 144062
rect 178309 144059 178375 144062
rect 22737 142898 22803 142901
rect 178401 142898 178467 142901
rect 22737 142896 178467 142898
rect 22737 142840 22742 142896
rect 22798 142840 178406 142896
rect 178462 142840 178467 142896
rect 22737 142838 178467 142840
rect 22737 142835 22803 142838
rect 178401 142835 178467 142838
rect 113909 142762 113975 142765
rect 439497 142762 439563 142765
rect 113909 142760 439563 142762
rect 113909 142704 113914 142760
rect 113970 142704 439502 142760
rect 439558 142704 439563 142760
rect 113909 142702 439563 142704
rect 113909 142699 113975 142702
rect 439497 142699 439563 142702
rect 351913 142218 351979 142221
rect 355685 142218 355751 142221
rect 351913 142216 355751 142218
rect 351913 142160 351918 142216
rect 351974 142160 355690 142216
rect 355746 142160 355751 142216
rect 351913 142158 355751 142160
rect 351913 142155 351979 142158
rect 355685 142155 355751 142158
rect 40493 141538 40559 141541
rect 176929 141538 176995 141541
rect 40493 141536 176995 141538
rect 40493 141480 40498 141536
rect 40554 141480 176934 141536
rect 176990 141480 176995 141536
rect 40493 141478 176995 141480
rect 40493 141475 40559 141478
rect 176929 141475 176995 141478
rect 115473 141402 115539 141405
rect 543457 141402 543523 141405
rect 115473 141400 543523 141402
rect 115473 141344 115478 141400
rect 115534 141344 543462 141400
rect 543518 141344 543523 141400
rect 115473 141342 543523 141344
rect 115473 141339 115539 141342
rect 543457 141339 543523 141342
rect 70761 140858 70827 140861
rect 73153 140858 73219 140861
rect 70761 140856 73219 140858
rect 70761 140800 70766 140856
rect 70822 140800 73158 140856
rect 73214 140800 73219 140856
rect 70761 140798 73219 140800
rect 70761 140795 70827 140798
rect 73153 140795 73219 140798
rect 116669 139362 116735 139365
rect 583520 139362 584960 139452
rect 116669 139360 584960 139362
rect 116669 139304 116674 139360
rect 116730 139304 584960 139360
rect 116669 139302 584960 139304
rect 116669 139299 116735 139302
rect 583520 139212 584960 139302
rect 18597 138682 18663 138685
rect 178585 138682 178651 138685
rect 18597 138680 178651 138682
rect 18597 138624 18602 138680
rect 18658 138624 178590 138680
rect 178646 138624 178651 138680
rect 18597 138622 178651 138624
rect 18597 138619 18663 138622
rect 178585 138619 178651 138622
rect 349153 138138 349219 138141
rect 351913 138138 351979 138141
rect 349153 138136 351979 138138
rect 349153 138080 349158 138136
rect 349214 138080 351918 138136
rect 351974 138080 351979 138136
rect 349153 138078 351979 138080
rect 349153 138075 349219 138078
rect 351913 138075 351979 138078
rect 125593 137594 125659 137597
rect 135846 137594 135852 137596
rect 125593 137592 135852 137594
rect 125593 137536 125598 137592
rect 125654 137536 135852 137592
rect 125593 137534 135852 137536
rect 125593 137531 125659 137534
rect 135846 137532 135852 137534
rect 135916 137532 135922 137596
rect 122465 137458 122531 137461
rect 136030 137458 136036 137460
rect 122465 137456 136036 137458
rect 122465 137400 122470 137456
rect 122526 137400 136036 137456
rect 122465 137398 136036 137400
rect 122465 137395 122531 137398
rect 136030 137396 136036 137398
rect 136100 137396 136106 137460
rect 141918 137396 141924 137460
rect 141988 137458 141994 137460
rect 167821 137458 167887 137461
rect 141988 137456 167887 137458
rect 141988 137400 167826 137456
rect 167882 137400 167887 137456
rect 141988 137398 167887 137400
rect 141988 137396 141994 137398
rect 167821 137395 167887 137398
rect 113725 137322 113791 137325
rect 446397 137322 446463 137325
rect 113725 137320 446463 137322
rect 113725 137264 113730 137320
rect 113786 137264 446402 137320
rect 446458 137264 446463 137320
rect 113725 137262 446463 137264
rect 113725 137259 113791 137262
rect 446397 137259 446463 137262
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 15837 136234 15903 136237
rect 178493 136234 178559 136237
rect 15837 136232 178559 136234
rect 15837 136176 15842 136232
rect 15898 136176 178498 136232
rect 178554 136176 178559 136232
rect 15837 136174 178559 136176
rect 15837 136171 15903 136174
rect 178493 136171 178559 136174
rect 115381 136098 115447 136101
rect 413645 136098 413711 136101
rect 115381 136096 413711 136098
rect 115381 136040 115386 136096
rect 115442 136040 413650 136096
rect 413706 136040 413711 136096
rect 115381 136038 413711 136040
rect 115381 136035 115447 136038
rect 413645 136035 413711 136038
rect 115565 135962 115631 135965
rect 580625 135962 580691 135965
rect 115565 135960 580691 135962
rect 115565 135904 115570 135960
rect 115626 135904 580630 135960
rect 580686 135904 580691 135960
rect 115565 135902 580691 135904
rect 115565 135899 115631 135902
rect 580625 135899 580691 135902
rect 345657 135146 345723 135149
rect 349061 135146 349127 135149
rect 345657 135144 349127 135146
rect 345657 135088 345662 135144
rect 345718 135088 349066 135144
rect 349122 135088 349127 135144
rect 345657 135086 349127 135088
rect 345657 135083 345723 135086
rect 349061 135083 349127 135086
rect 73153 134466 73219 134469
rect 176653 134466 176719 134469
rect 73153 134464 176719 134466
rect 73153 134408 73158 134464
rect 73214 134408 176658 134464
rect 176714 134408 176719 134464
rect 73153 134406 176719 134408
rect 73153 134403 73219 134406
rect 176653 134403 176719 134406
rect 15837 134330 15903 134333
rect 178033 134330 178099 134333
rect 15837 134328 178099 134330
rect 15837 134272 15842 134328
rect 15898 134272 178038 134328
rect 178094 134272 178099 134328
rect 15837 134270 178099 134272
rect 15837 134267 15903 134270
rect 178033 134267 178099 134270
rect 113817 133242 113883 133245
rect 113817 133240 116226 133242
rect 113817 133184 113822 133240
rect 113878 133184 116226 133240
rect 113817 133182 116226 133184
rect 113817 133179 113883 133182
rect 3601 133106 3667 133109
rect 17953 133106 18019 133109
rect 3601 133104 18019 133106
rect 3601 133048 3606 133104
rect 3662 133048 17958 133104
rect 18014 133048 18019 133104
rect 3601 133046 18019 133048
rect 3601 133043 3667 133046
rect 17953 133043 18019 133046
rect 116166 132600 116226 133182
rect 175782 132562 175842 132600
rect 177021 132562 177087 132565
rect 175782 132560 177087 132562
rect 175782 132504 177026 132560
rect 177082 132504 177087 132560
rect 175782 132502 177087 132504
rect 177021 132499 177087 132502
rect 3601 131202 3667 131205
rect 178953 131202 179019 131205
rect 3601 131200 116226 131202
rect 3601 131144 3606 131200
rect 3662 131144 116226 131200
rect 3601 131142 116226 131144
rect 3601 131139 3667 131142
rect 116166 131104 116226 131142
rect 175782 131200 179019 131202
rect 175782 131144 178958 131200
rect 179014 131144 179019 131200
rect 175782 131142 179019 131144
rect 175782 131104 175842 131142
rect 178953 131139 179019 131142
rect 113817 129842 113883 129845
rect 116485 129842 116551 129845
rect 113817 129840 116551 129842
rect 113817 129784 113822 129840
rect 113878 129784 116490 129840
rect 116546 129784 116551 129840
rect 113817 129782 116551 129784
rect 113817 129779 113883 129782
rect 116485 129779 116551 129782
rect 178033 129706 178099 129709
rect 175782 129704 178099 129706
rect 175782 129648 178038 129704
rect 178094 129648 178099 129704
rect 175782 129646 178099 129648
rect 175782 129608 175842 129646
rect 178033 129643 178099 129646
rect 3693 128482 3759 128485
rect 116166 128482 116226 129608
rect 3693 128480 116226 128482
rect 3693 128424 3698 128480
rect 3754 128424 116226 128480
rect 3693 128422 116226 128424
rect 3693 128419 3759 128422
rect 176745 128346 176811 128349
rect 175782 128344 176811 128346
rect 175782 128288 176750 128344
rect 176806 128288 176811 128344
rect 175782 128286 176811 128288
rect 175782 128112 175842 128286
rect 176745 128283 176811 128286
rect 3785 127122 3851 127125
rect 116166 127122 116226 128112
rect 3785 127120 116226 127122
rect 3785 127064 3790 127120
rect 3846 127064 116226 127120
rect 3785 127062 116226 127064
rect 3785 127059 3851 127062
rect 17953 126986 18019 126989
rect 175365 126986 175431 126989
rect 17953 126984 116226 126986
rect 17953 126928 17958 126984
rect 18014 126928 116226 126984
rect 17953 126926 116226 126928
rect 17953 126923 18019 126926
rect 116166 126616 116226 126926
rect 175365 126984 175474 126986
rect 175365 126928 175370 126984
rect 175426 126928 175474 126984
rect 175365 126923 175474 126928
rect 175414 126616 175474 126923
rect 184197 126034 184263 126037
rect 583520 126034 584960 126124
rect 184197 126032 584960 126034
rect 184197 125976 184202 126032
rect 184258 125976 584960 126032
rect 184197 125974 584960 125976
rect 184197 125971 184263 125974
rect 583520 125884 584960 125974
rect 46197 125490 46263 125493
rect 176837 125490 176903 125493
rect 46197 125488 116226 125490
rect 46197 125432 46202 125488
rect 46258 125432 116226 125488
rect 46197 125430 116226 125432
rect 46197 125427 46263 125430
rect 116166 125120 116226 125430
rect 175782 125488 176903 125490
rect 175782 125432 176842 125488
rect 176898 125432 176903 125488
rect 175782 125430 176903 125432
rect 175782 125120 175842 125430
rect 176837 125427 176903 125430
rect 22829 124130 22895 124133
rect 178769 124130 178835 124133
rect 22829 124128 116226 124130
rect 22829 124072 22834 124128
rect 22890 124072 116226 124128
rect 22829 124070 116226 124072
rect 22829 124067 22895 124070
rect -960 123572 480 123812
rect 116166 123624 116226 124070
rect 175782 124128 178835 124130
rect 175782 124072 178774 124128
rect 178830 124072 178835 124128
rect 175782 124070 178835 124072
rect 175782 123624 175842 124070
rect 178769 124067 178835 124070
rect 31109 122770 31175 122773
rect 31109 122768 116226 122770
rect 31109 122712 31114 122768
rect 31170 122712 116226 122768
rect 31109 122710 116226 122712
rect 31109 122707 31175 122710
rect 116166 122128 116226 122710
rect 178677 122498 178743 122501
rect 175782 122496 178743 122498
rect 175782 122440 178682 122496
rect 178738 122440 178743 122496
rect 175782 122438 178743 122440
rect 175782 122128 175842 122438
rect 178677 122435 178743 122438
rect 14457 121410 14523 121413
rect 14457 121408 116226 121410
rect 14457 121352 14462 121408
rect 14518 121352 116226 121408
rect 14457 121350 116226 121352
rect 14457 121347 14523 121350
rect 116166 120632 116226 121350
rect 177849 121274 177915 121277
rect 175782 121272 177915 121274
rect 175782 121216 177854 121272
rect 177910 121216 177915 121272
rect 175782 121214 177915 121216
rect 175782 120632 175842 121214
rect 177849 121211 177915 121214
rect 11697 120050 11763 120053
rect 11697 120048 116226 120050
rect 11697 119992 11702 120048
rect 11758 119992 116226 120048
rect 11697 119990 116226 119992
rect 11697 119987 11763 119990
rect 116166 119136 116226 119990
rect 178217 119778 178283 119781
rect 175782 119776 178283 119778
rect 175782 119720 178222 119776
rect 178278 119720 178283 119776
rect 175782 119718 178283 119720
rect 175782 119136 175842 119718
rect 178217 119715 178283 119718
rect 175917 118826 175983 118829
rect 178217 118826 178283 118829
rect 175917 118824 178283 118826
rect 175917 118768 175922 118824
rect 175978 118768 178222 118824
rect 178278 118768 178283 118824
rect 175917 118766 178283 118768
rect 175917 118763 175983 118766
rect 178217 118763 178283 118766
rect 4981 118690 5047 118693
rect 4981 118688 116226 118690
rect 4981 118632 4986 118688
rect 5042 118632 116226 118688
rect 4981 118630 116226 118632
rect 4981 118627 5047 118630
rect 116166 117640 116226 118630
rect 178309 118282 178375 118285
rect 175782 118280 178375 118282
rect 175782 118224 178314 118280
rect 178370 118224 178375 118280
rect 175782 118222 178375 118224
rect 175782 117640 175842 118222
rect 178309 118219 178375 118222
rect 4797 117194 4863 117197
rect 4797 117192 116226 117194
rect 4797 117136 4802 117192
rect 4858 117136 116226 117192
rect 4797 117134 116226 117136
rect 4797 117131 4863 117134
rect 116166 116144 116226 117134
rect 178401 116786 178467 116789
rect 175782 116784 178467 116786
rect 175782 116728 178406 116784
rect 178462 116728 178467 116784
rect 175782 116726 178467 116728
rect 175782 116144 175842 116726
rect 178401 116723 178467 116726
rect 337377 116514 337443 116517
rect 345657 116514 345723 116517
rect 337377 116512 345723 116514
rect 337377 116456 337382 116512
rect 337438 116456 345662 116512
rect 345718 116456 345723 116512
rect 337377 116454 345723 116456
rect 337377 116451 337443 116454
rect 345657 116451 345723 116454
rect 25589 115834 25655 115837
rect 25589 115832 116226 115834
rect 25589 115776 25594 115832
rect 25650 115776 116226 115832
rect 25589 115774 116226 115776
rect 25589 115771 25655 115774
rect 116166 114648 116226 115774
rect 178585 115290 178651 115293
rect 175782 115288 178651 115290
rect 175782 115232 178590 115288
rect 178646 115232 178651 115288
rect 175782 115230 178651 115232
rect 175782 114648 175842 115230
rect 178585 115227 178651 115230
rect 29637 113114 29703 113117
rect 116166 113114 116226 113152
rect 29637 113112 116226 113114
rect 29637 113056 29642 113112
rect 29698 113056 116226 113112
rect 29637 113054 116226 113056
rect 175782 113114 175842 113152
rect 178493 113114 178559 113117
rect 175782 113112 178559 113114
rect 175782 113056 178498 113112
rect 178554 113056 178559 113112
rect 175782 113054 178559 113056
rect 29637 113051 29703 113054
rect 178493 113051 178559 113054
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect 26877 111754 26943 111757
rect 176929 111754 176995 111757
rect 26877 111752 116226 111754
rect 26877 111696 26882 111752
rect 26938 111696 116226 111752
rect 26877 111694 116226 111696
rect 26877 111691 26943 111694
rect 116166 111656 116226 111694
rect 175782 111752 176995 111754
rect 175782 111696 176934 111752
rect 176990 111696 176995 111752
rect 175782 111694 176995 111696
rect 175782 111656 175842 111694
rect 176929 111691 176995 111694
rect -960 110666 480 110756
rect 15837 110666 15903 110669
rect -960 110664 15903 110666
rect -960 110608 15842 110664
rect 15898 110608 15903 110664
rect -960 110606 15903 110608
rect -960 110516 480 110606
rect 15837 110603 15903 110606
rect 24301 110394 24367 110397
rect 178125 110394 178191 110397
rect 24301 110392 116226 110394
rect 24301 110336 24306 110392
rect 24362 110336 116226 110392
rect 24301 110334 116226 110336
rect 24301 110331 24367 110334
rect 116166 110160 116226 110334
rect 175782 110392 178191 110394
rect 175782 110336 178130 110392
rect 178186 110336 178191 110392
rect 175782 110334 178191 110336
rect 175782 110160 175842 110334
rect 178125 110331 178191 110334
rect 45093 109034 45159 109037
rect 178217 109034 178283 109037
rect 45093 109032 116226 109034
rect 45093 108976 45098 109032
rect 45154 108976 116226 109032
rect 45093 108974 116226 108976
rect 45093 108971 45159 108974
rect 116166 108664 116226 108974
rect 175782 109032 178283 109034
rect 175782 108976 178222 109032
rect 178278 108976 178283 109032
rect 175782 108974 178283 108976
rect 175782 108664 175842 108974
rect 178217 108971 178283 108974
rect 331213 109034 331279 109037
rect 337377 109034 337443 109037
rect 331213 109032 337443 109034
rect 331213 108976 331218 109032
rect 331274 108976 337382 109032
rect 337438 108976 337443 109032
rect 331213 108974 337443 108976
rect 331213 108971 331279 108974
rect 337377 108971 337443 108974
rect 45369 107538 45435 107541
rect 176653 107538 176719 107541
rect 45369 107536 116226 107538
rect 45369 107480 45374 107536
rect 45430 107480 116226 107536
rect 45369 107478 116226 107480
rect 45369 107475 45435 107478
rect 116166 107168 116226 107478
rect 175782 107536 176719 107538
rect 175782 107480 176658 107536
rect 176714 107480 176719 107536
rect 175782 107478 176719 107480
rect 175782 107168 175842 107478
rect 176653 107475 176719 107478
rect 322933 106858 322999 106861
rect 331213 106858 331279 106861
rect 322933 106856 331279 106858
rect 322933 106800 322938 106856
rect 322994 106800 331218 106856
rect 331274 106800 331279 106856
rect 322933 106798 331279 106800
rect 322933 106795 322999 106798
rect 331213 106795 331279 106798
rect 44909 106178 44975 106181
rect 322933 106178 322999 106181
rect 44909 106176 116226 106178
rect 44909 106120 44914 106176
rect 44970 106120 116226 106176
rect 44909 106118 116226 106120
rect 44909 106115 44975 106118
rect 116166 105672 116226 106118
rect 175782 106176 322999 106178
rect 175782 106120 322938 106176
rect 322994 106120 322999 106176
rect 175782 106118 322999 106120
rect 175782 105672 175842 106118
rect 322933 106115 322999 106118
rect 45737 104818 45803 104821
rect 396533 104818 396599 104821
rect 45737 104816 116226 104818
rect 45737 104760 45742 104816
rect 45798 104760 116226 104816
rect 45737 104758 116226 104760
rect 45737 104755 45803 104758
rect 116166 104176 116226 104758
rect 175782 104816 396599 104818
rect 175782 104760 396538 104816
rect 396594 104760 396599 104816
rect 175782 104758 396599 104760
rect 175782 104176 175842 104758
rect 396533 104755 396599 104758
rect 416037 103458 416103 103461
rect 175782 103456 416103 103458
rect 175782 103400 416042 103456
rect 416098 103400 416103 103456
rect 175782 103398 416103 103400
rect 114369 103186 114435 103189
rect 114369 103184 116226 103186
rect 114369 103128 114374 103184
rect 114430 103128 116226 103184
rect 114369 103126 116226 103128
rect 114369 103123 114435 103126
rect 116166 102680 116226 103126
rect 175782 102680 175842 103398
rect 416037 103395 416103 103398
rect 414657 102098 414723 102101
rect 180750 102096 414723 102098
rect 180750 102040 414662 102096
rect 414718 102040 414723 102096
rect 180750 102038 414723 102040
rect 180750 101962 180810 102038
rect 414657 102035 414723 102038
rect 175782 101902 180810 101962
rect 115381 101826 115447 101829
rect 115381 101824 116226 101826
rect 115381 101768 115386 101824
rect 115442 101768 116226 101824
rect 115381 101766 116226 101768
rect 115381 101763 115447 101766
rect 116166 101184 116226 101766
rect 175782 101184 175842 101902
rect 406377 100738 406443 100741
rect 180750 100736 406443 100738
rect 180750 100680 406382 100736
rect 406438 100680 406443 100736
rect 180750 100678 406443 100680
rect 180750 100466 180810 100678
rect 406377 100675 406443 100678
rect 175782 100406 180810 100466
rect 116485 100330 116551 100333
rect 116485 100328 116594 100330
rect 116485 100272 116490 100328
rect 116546 100272 116594 100328
rect 116485 100267 116594 100272
rect 116534 99688 116594 100267
rect 175782 99688 175842 100406
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 544377 99378 544443 99381
rect 180750 99376 544443 99378
rect 180750 99320 544382 99376
rect 544438 99320 544443 99376
rect 583520 99364 584960 99454
rect 180750 99318 544443 99320
rect 180750 98970 180810 99318
rect 544377 99315 544443 99318
rect 175782 98910 180810 98970
rect 115473 98834 115539 98837
rect 115473 98832 116226 98834
rect 115473 98776 115478 98832
rect 115534 98776 116226 98832
rect 115473 98774 116226 98776
rect 115473 98771 115539 98774
rect 116166 98192 116226 98774
rect 175782 98192 175842 98910
rect 404997 97882 405063 97885
rect 180750 97880 405063 97882
rect 180750 97824 405002 97880
rect 405058 97824 405063 97880
rect 180750 97822 405063 97824
rect -960 97610 480 97700
rect 3785 97610 3851 97613
rect -960 97608 3851 97610
rect -960 97552 3790 97608
rect 3846 97552 3851 97608
rect -960 97550 3851 97552
rect -960 97460 480 97550
rect 3785 97547 3851 97550
rect 180750 97474 180810 97822
rect 404997 97819 405063 97822
rect 175782 97414 180810 97474
rect 115749 96726 115815 96729
rect 115749 96724 116196 96726
rect 115749 96668 115754 96724
rect 115810 96668 116196 96724
rect 175782 96696 175842 97414
rect 115749 96666 116196 96668
rect 115749 96663 115815 96666
rect 115657 95230 115723 95233
rect 115657 95228 116196 95230
rect 115657 95172 115662 95228
rect 115718 95172 116196 95228
rect 115657 95170 116196 95172
rect 115657 95167 115723 95170
rect 175782 95162 175842 95200
rect 403617 95162 403683 95165
rect 175782 95160 403683 95162
rect 175782 95104 403622 95160
rect 403678 95104 403683 95160
rect 175782 95102 403683 95104
rect 403617 95099 403683 95102
rect 400857 93802 400923 93805
rect 175782 93800 400923 93802
rect 175782 93744 400862 93800
rect 400918 93744 400923 93800
rect 175782 93742 400923 93744
rect 115841 93734 115907 93737
rect 115841 93732 116196 93734
rect 115841 93676 115846 93732
rect 115902 93676 116196 93732
rect 175782 93704 175842 93742
rect 400857 93739 400923 93742
rect 115841 93674 116196 93676
rect 115841 93671 115907 93674
rect 115565 92442 115631 92445
rect 399477 92442 399543 92445
rect 115565 92440 116226 92442
rect 115565 92384 115570 92440
rect 115626 92384 116226 92440
rect 115565 92382 116226 92384
rect 115565 92379 115631 92382
rect 116166 92208 116226 92382
rect 175782 92440 399543 92442
rect 175782 92384 399482 92440
rect 399538 92384 399543 92440
rect 175782 92382 399543 92384
rect 175782 92208 175842 92382
rect 399477 92379 399543 92382
rect 113725 91082 113791 91085
rect 411897 91082 411963 91085
rect 113725 91080 116226 91082
rect 113725 91024 113730 91080
rect 113786 91024 116226 91080
rect 113725 91022 116226 91024
rect 113725 91019 113791 91022
rect 116166 90712 116226 91022
rect 175782 91080 411963 91082
rect 175782 91024 411902 91080
rect 411958 91024 411963 91080
rect 175782 91022 411963 91024
rect 175782 90712 175842 91022
rect 411897 91019 411963 91022
rect 113909 89722 113975 89725
rect 420177 89722 420243 89725
rect 113909 89720 116226 89722
rect 113909 89664 113914 89720
rect 113970 89664 116226 89720
rect 113909 89662 116226 89664
rect 113909 89659 113975 89662
rect 116166 89216 116226 89662
rect 175782 89720 420243 89722
rect 175782 89664 420182 89720
rect 420238 89664 420243 89720
rect 175782 89662 420243 89664
rect 175782 89216 175842 89662
rect 420177 89659 420243 89662
rect 114001 88226 114067 88229
rect 409137 88226 409203 88229
rect 114001 88224 116226 88226
rect 114001 88168 114006 88224
rect 114062 88168 116226 88224
rect 114001 88166 116226 88168
rect 114001 88163 114067 88166
rect 116166 87720 116226 88166
rect 175782 88224 409203 88226
rect 175782 88168 409142 88224
rect 409198 88168 409203 88224
rect 175782 88166 409203 88168
rect 175782 87720 175842 88166
rect 409137 88163 409203 88166
rect 114093 86866 114159 86869
rect 407757 86866 407823 86869
rect 114093 86864 116226 86866
rect 114093 86808 114098 86864
rect 114154 86808 116226 86864
rect 114093 86806 116226 86808
rect 114093 86803 114159 86806
rect 116166 86224 116226 86806
rect 175782 86864 407823 86866
rect 175782 86808 407762 86864
rect 407818 86808 407823 86864
rect 175782 86806 407823 86808
rect 175782 86224 175842 86806
rect 407757 86803 407823 86806
rect 178493 86186 178559 86189
rect 583520 86186 584960 86276
rect 178493 86184 584960 86186
rect 178493 86128 178498 86184
rect 178554 86128 584960 86184
rect 178493 86126 584960 86128
rect 178493 86123 178559 86126
rect 583520 86036 584960 86126
rect 188337 85506 188403 85509
rect 175782 85504 188403 85506
rect 175782 85448 188342 85504
rect 188398 85448 188403 85504
rect 175782 85446 188403 85448
rect 114185 85370 114251 85373
rect 114185 85368 116226 85370
rect 114185 85312 114190 85368
rect 114246 85312 116226 85368
rect 114185 85310 116226 85312
rect 114185 85307 114251 85310
rect -960 84690 480 84780
rect 116166 84728 116226 85310
rect 175782 84728 175842 85446
rect 188337 85443 188403 85446
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 185577 84010 185643 84013
rect 175782 84008 185643 84010
rect 175782 83952 185582 84008
rect 185638 83952 185643 84008
rect 175782 83950 185643 83952
rect 114461 83738 114527 83741
rect 114461 83736 116226 83738
rect 114461 83680 114466 83736
rect 114522 83680 116226 83736
rect 114461 83678 116226 83680
rect 114461 83675 114527 83678
rect 116166 83232 116226 83678
rect 175782 83232 175842 83950
rect 185577 83947 185643 83950
rect 184197 82514 184263 82517
rect 175782 82512 184263 82514
rect 175782 82456 184202 82512
rect 184258 82456 184263 82512
rect 175782 82454 184263 82456
rect 114277 82378 114343 82381
rect 114277 82376 116226 82378
rect 114277 82320 114282 82376
rect 114338 82320 116226 82376
rect 114277 82318 116226 82320
rect 114277 82315 114343 82318
rect 116166 81736 116226 82318
rect 175782 81736 175842 82454
rect 184197 82451 184263 82454
rect 113817 80882 113883 80885
rect 178493 80882 178559 80885
rect 113817 80880 116226 80882
rect 113817 80824 113822 80880
rect 113878 80824 116226 80880
rect 113817 80822 116226 80824
rect 113817 80819 113883 80822
rect 116166 80240 116226 80822
rect 175782 80880 178559 80882
rect 175782 80824 178498 80880
rect 178554 80824 178559 80880
rect 175782 80822 178559 80824
rect 175782 80240 175842 80822
rect 178493 80819 178559 80822
rect 116534 78165 116594 78744
rect 175782 78706 175842 78744
rect 178769 78706 178835 78709
rect 175782 78704 178835 78706
rect 175782 78648 178774 78704
rect 178830 78648 178835 78704
rect 175782 78646 178835 78648
rect 178769 78643 178835 78646
rect 116485 78160 116594 78165
rect 116485 78104 116490 78160
rect 116546 78104 116594 78160
rect 116485 78102 116594 78104
rect 116485 78099 116551 78102
rect 114369 76666 114435 76669
rect 116166 76666 116226 77248
rect 114369 76664 116226 76666
rect 114369 76608 114374 76664
rect 114430 76608 116226 76664
rect 114369 76606 116226 76608
rect 175782 76666 175842 77248
rect 178861 76666 178927 76669
rect 175782 76664 178927 76666
rect 175782 76608 178866 76664
rect 178922 76608 178927 76664
rect 175782 76606 178927 76608
rect 114369 76603 114435 76606
rect 178861 76603 178927 76606
rect 114461 75170 114527 75173
rect 116166 75170 116226 75752
rect 116485 75578 116551 75581
rect 170673 75578 170739 75581
rect 116485 75576 170739 75578
rect 116485 75520 116490 75576
rect 116546 75520 170678 75576
rect 170734 75520 170739 75576
rect 116485 75518 170739 75520
rect 116485 75515 116551 75518
rect 170673 75515 170739 75518
rect 169334 75380 169340 75444
rect 169404 75442 169410 75444
rect 170673 75442 170739 75445
rect 169404 75440 170739 75442
rect 169404 75384 170678 75440
rect 170734 75384 170739 75440
rect 169404 75382 170739 75384
rect 169404 75380 169410 75382
rect 170673 75379 170739 75382
rect 147438 75244 147444 75308
rect 147508 75306 147514 75308
rect 228725 75306 228791 75309
rect 147508 75304 228791 75306
rect 147508 75248 228730 75304
rect 228786 75248 228791 75304
rect 147508 75246 228791 75248
rect 147508 75244 147514 75246
rect 228725 75243 228791 75246
rect 114461 75168 116226 75170
rect 114461 75112 114466 75168
rect 114522 75112 116226 75168
rect 114461 75110 116226 75112
rect 114461 75107 114527 75110
rect 160870 75108 160876 75172
rect 160940 75170 160946 75172
rect 196801 75170 196867 75173
rect 160940 75168 196867 75170
rect 160940 75112 196806 75168
rect 196862 75112 196867 75168
rect 160940 75110 196867 75112
rect 160940 75108 160946 75110
rect 196801 75107 196867 75110
rect 179045 75034 179111 75037
rect 137970 75032 179111 75034
rect 137970 74976 179050 75032
rect 179106 74976 179111 75032
rect 137970 74974 179111 74976
rect 135437 74898 135503 74901
rect 137970 74898 138030 74974
rect 179045 74971 179111 74974
rect 135437 74896 138030 74898
rect 135437 74840 135442 74896
rect 135498 74840 138030 74896
rect 135437 74838 138030 74840
rect 157701 74898 157767 74901
rect 158846 74898 158852 74900
rect 157701 74896 158852 74898
rect 157701 74840 157706 74896
rect 157762 74840 158852 74896
rect 157701 74838 158852 74840
rect 135437 74835 135503 74838
rect 157701 74835 157767 74838
rect 158846 74836 158852 74838
rect 158916 74836 158922 74900
rect 161422 74836 161428 74900
rect 161492 74898 161498 74900
rect 214465 74898 214531 74901
rect 161492 74896 214531 74898
rect 161492 74840 214470 74896
rect 214526 74840 214531 74896
rect 161492 74838 214531 74840
rect 161492 74836 161498 74838
rect 214465 74835 214531 74838
rect 155902 74700 155908 74764
rect 155972 74762 155978 74764
rect 218053 74762 218119 74765
rect 155972 74760 218119 74762
rect 155972 74704 218058 74760
rect 218114 74704 218119 74760
rect 155972 74702 218119 74704
rect 155972 74700 155978 74702
rect 218053 74699 218119 74702
rect 152273 74626 152339 74629
rect 157190 74626 157196 74628
rect 152273 74624 157196 74626
rect 152273 74568 152278 74624
rect 152334 74568 157196 74624
rect 152273 74566 157196 74568
rect 152273 74563 152339 74566
rect 157190 74564 157196 74566
rect 157260 74564 157266 74628
rect 167545 74626 167611 74629
rect 169334 74626 169340 74628
rect 167545 74624 169340 74626
rect 167545 74568 167550 74624
rect 167606 74568 169340 74624
rect 167545 74566 169340 74568
rect 167545 74563 167611 74566
rect 169334 74564 169340 74566
rect 169404 74564 169410 74628
rect 169477 74626 169543 74629
rect 170397 74626 170463 74629
rect 169477 74624 170463 74626
rect 169477 74568 169482 74624
rect 169538 74568 170402 74624
rect 170458 74568 170463 74624
rect 169477 74566 170463 74568
rect 169477 74563 169543 74566
rect 170397 74563 170463 74566
rect 21357 74490 21423 74493
rect 169845 74490 169911 74493
rect 21357 74488 169911 74490
rect 21357 74432 21362 74488
rect 21418 74432 169850 74488
rect 169906 74432 169911 74488
rect 21357 74430 169911 74432
rect 21357 74427 21423 74430
rect 169845 74427 169911 74430
rect 134977 74354 135043 74357
rect 173157 74354 173223 74357
rect 134977 74352 173223 74354
rect 134977 74296 134982 74352
rect 135038 74296 173162 74352
rect 173218 74296 173223 74352
rect 134977 74294 173223 74296
rect 134977 74291 135043 74294
rect 173157 74291 173223 74294
rect 139577 74218 139643 74221
rect 232221 74218 232287 74221
rect 139577 74216 232287 74218
rect 139577 74160 139582 74216
rect 139638 74160 232226 74216
rect 232282 74160 232287 74216
rect 139577 74158 232287 74160
rect 139577 74155 139643 74158
rect 232221 74155 232287 74158
rect 142337 74082 142403 74085
rect 267733 74082 267799 74085
rect 142337 74080 267799 74082
rect 142337 74024 142342 74080
rect 142398 74024 267738 74080
rect 267794 74024 267799 74080
rect 142337 74022 267799 74024
rect 142337 74019 142403 74022
rect 267733 74019 267799 74022
rect 151486 73884 151492 73948
rect 151556 73946 151562 73948
rect 151629 73946 151695 73949
rect 151556 73944 151695 73946
rect 151556 73888 151634 73944
rect 151690 73888 151695 73944
rect 151556 73886 151695 73888
rect 151556 73884 151562 73886
rect 151629 73883 151695 73886
rect 157190 73884 157196 73948
rect 157260 73946 157266 73948
rect 395337 73946 395403 73949
rect 157260 73944 395403 73946
rect 157260 73888 395342 73944
rect 395398 73888 395403 73944
rect 157260 73886 395403 73888
rect 157260 73884 157266 73886
rect 395337 73883 395403 73886
rect 158897 73810 158963 73813
rect 480529 73810 480595 73813
rect 158897 73808 480595 73810
rect 158897 73752 158902 73808
rect 158958 73752 480534 73808
rect 480590 73752 480595 73808
rect 158897 73750 480595 73752
rect 158897 73747 158963 73750
rect 480529 73747 480595 73750
rect 140262 73612 140268 73676
rect 140332 73674 140338 73676
rect 140681 73674 140747 73677
rect 140332 73672 140747 73674
rect 140332 73616 140686 73672
rect 140742 73616 140747 73672
rect 140332 73614 140747 73616
rect 140332 73612 140338 73614
rect 140681 73611 140747 73614
rect 123661 73540 123727 73541
rect 139117 73540 139183 73541
rect 140497 73540 140563 73541
rect 123661 73536 123708 73540
rect 123772 73538 123778 73540
rect 123661 73480 123666 73536
rect 123661 73476 123708 73480
rect 123772 73478 123818 73538
rect 139117 73536 139164 73540
rect 139228 73538 139234 73540
rect 140446 73538 140452 73540
rect 139117 73480 139122 73536
rect 123772 73476 123778 73478
rect 139117 73476 139164 73480
rect 139228 73478 139274 73538
rect 140406 73478 140452 73538
rect 140516 73536 140563 73540
rect 140558 73480 140563 73536
rect 139228 73476 139234 73478
rect 140446 73476 140452 73478
rect 140516 73476 140563 73480
rect 141182 73476 141188 73540
rect 141252 73538 141258 73540
rect 142061 73538 142127 73541
rect 141252 73536 142127 73538
rect 141252 73480 142066 73536
rect 142122 73480 142127 73536
rect 141252 73478 142127 73480
rect 141252 73476 141258 73478
rect 123661 73475 123727 73476
rect 139117 73475 139183 73476
rect 140497 73475 140563 73476
rect 142061 73475 142127 73478
rect 153101 73538 153167 73541
rect 161197 73538 161263 73541
rect 161606 73538 161612 73540
rect 153101 73536 160110 73538
rect 153101 73480 153106 73536
rect 153162 73480 160110 73536
rect 153101 73478 160110 73480
rect 153101 73475 153167 73478
rect 139209 73402 139275 73405
rect 139342 73402 139348 73404
rect 139209 73400 139348 73402
rect 139209 73344 139214 73400
rect 139270 73344 139348 73400
rect 139209 73342 139348 73344
rect 139209 73339 139275 73342
rect 139342 73340 139348 73342
rect 139412 73340 139418 73404
rect 140078 73340 140084 73404
rect 140148 73402 140154 73404
rect 140405 73402 140471 73405
rect 140148 73400 140471 73402
rect 140148 73344 140410 73400
rect 140466 73344 140471 73400
rect 140148 73342 140471 73344
rect 140148 73340 140154 73342
rect 140405 73339 140471 73342
rect 140589 73404 140655 73405
rect 158897 73404 158963 73405
rect 140589 73400 140636 73404
rect 140700 73402 140706 73404
rect 140589 73344 140594 73400
rect 140589 73340 140636 73344
rect 140700 73342 140746 73402
rect 140700 73340 140706 73342
rect 158846 73340 158852 73404
rect 158916 73402 158963 73404
rect 160050 73402 160110 73478
rect 161197 73536 161612 73538
rect 161197 73480 161202 73536
rect 161258 73480 161612 73536
rect 161197 73478 161612 73480
rect 161197 73475 161263 73478
rect 161606 73476 161612 73478
rect 161676 73476 161682 73540
rect 166206 73476 166212 73540
rect 166276 73538 166282 73540
rect 166809 73538 166875 73541
rect 166276 73536 166875 73538
rect 166276 73480 166814 73536
rect 166870 73480 166875 73536
rect 166276 73478 166875 73480
rect 166276 73476 166282 73478
rect 166809 73475 166875 73478
rect 306741 73402 306807 73405
rect 158916 73400 159008 73402
rect 158958 73344 159008 73400
rect 158916 73342 159008 73344
rect 160050 73400 306807 73402
rect 160050 73344 306746 73400
rect 306802 73344 306807 73400
rect 160050 73342 306807 73344
rect 158916 73340 158963 73342
rect 140589 73339 140655 73340
rect 158897 73339 158963 73340
rect 306741 73339 306807 73342
rect 139853 73266 139919 73269
rect 157701 73266 157767 73269
rect 161289 73268 161355 73269
rect 161238 73266 161244 73268
rect 139853 73264 157767 73266
rect 139853 73208 139858 73264
rect 139914 73208 157706 73264
rect 157762 73208 157767 73264
rect 139853 73206 157767 73208
rect 161198 73206 161244 73266
rect 161308 73264 161355 73268
rect 161350 73208 161355 73264
rect 139853 73203 139919 73206
rect 157701 73203 157767 73206
rect 161238 73204 161244 73206
rect 161308 73204 161355 73208
rect 161289 73203 161355 73204
rect 161430 73206 164250 73266
rect 3417 73130 3483 73133
rect 117865 73130 117931 73133
rect 124305 73130 124371 73133
rect 3417 73128 117931 73130
rect 3417 73072 3422 73128
rect 3478 73072 117870 73128
rect 117926 73072 117931 73128
rect 3417 73070 117931 73072
rect 3417 73067 3483 73070
rect 117865 73067 117931 73070
rect 118006 73128 124371 73130
rect 118006 73072 124310 73128
rect 124366 73072 124371 73128
rect 118006 73070 124371 73072
rect 8109 72994 8175 72997
rect 118006 72994 118066 73070
rect 124305 73067 124371 73070
rect 129733 73130 129799 73133
rect 139301 73130 139367 73133
rect 147438 73130 147444 73132
rect 129733 73128 129842 73130
rect 129733 73072 129738 73128
rect 129794 73072 129842 73128
rect 129733 73067 129842 73072
rect 139301 73128 147444 73130
rect 139301 73072 139306 73128
rect 139362 73072 147444 73128
rect 139301 73070 147444 73072
rect 139301 73067 139367 73070
rect 147438 73068 147444 73070
rect 147508 73068 147514 73132
rect 147990 73068 147996 73132
rect 148060 73130 148066 73132
rect 148685 73130 148751 73133
rect 148060 73128 148751 73130
rect 148060 73072 148690 73128
rect 148746 73072 148751 73128
rect 148060 73070 148751 73072
rect 148060 73068 148066 73070
rect 148685 73067 148751 73070
rect 150433 73130 150499 73133
rect 157517 73132 157583 73133
rect 150433 73128 157442 73130
rect 150433 73072 150438 73128
rect 150494 73072 157442 73128
rect 150433 73070 157442 73072
rect 150433 73067 150499 73070
rect 8109 72992 118066 72994
rect 8109 72936 8114 72992
rect 8170 72936 118066 72992
rect 8109 72934 118066 72936
rect 120257 72994 120323 72997
rect 121913 72994 121979 72997
rect 126697 72994 126763 72997
rect 120257 72992 121979 72994
rect 120257 72936 120262 72992
rect 120318 72936 121918 72992
rect 121974 72936 121979 72992
rect 120257 72934 121979 72936
rect 8109 72931 8175 72934
rect 120257 72931 120323 72934
rect 121913 72931 121979 72934
rect 126654 72992 126763 72994
rect 126654 72936 126702 72992
rect 126758 72936 126763 72992
rect 126654 72931 126763 72936
rect 43437 72858 43503 72861
rect 123569 72858 123635 72861
rect 43437 72856 123635 72858
rect 43437 72800 43442 72856
rect 43498 72800 123574 72856
rect 123630 72800 123635 72856
rect 43437 72798 123635 72800
rect 43437 72795 43503 72798
rect 123569 72795 123635 72798
rect 124438 72796 124444 72860
rect 124508 72858 124514 72860
rect 124581 72858 124647 72861
rect 124508 72856 124647 72858
rect 124508 72800 124586 72856
rect 124642 72800 124647 72856
rect 124508 72798 124647 72800
rect 124508 72796 124514 72798
rect 124581 72795 124647 72798
rect 125542 72796 125548 72860
rect 125612 72858 125618 72860
rect 125685 72858 125751 72861
rect 125612 72856 125751 72858
rect 125612 72800 125690 72856
rect 125746 72800 125751 72856
rect 125612 72798 125751 72800
rect 125612 72796 125618 72798
rect 125685 72795 125751 72798
rect 120257 72722 120323 72725
rect 103470 72720 120323 72722
rect 103470 72664 120262 72720
rect 120318 72664 120323 72720
rect 103470 72662 120323 72664
rect 25497 72586 25563 72589
rect 103470 72586 103530 72662
rect 120257 72659 120323 72662
rect 121494 72660 121500 72724
rect 121564 72722 121570 72724
rect 121637 72722 121703 72725
rect 123201 72724 123267 72725
rect 123150 72722 123156 72724
rect 121564 72720 121703 72722
rect 121564 72664 121642 72720
rect 121698 72664 121703 72720
rect 121564 72662 121703 72664
rect 123110 72662 123156 72722
rect 123220 72720 123267 72724
rect 123262 72664 123267 72720
rect 121564 72660 121570 72662
rect 121637 72659 121703 72662
rect 123150 72660 123156 72662
rect 123220 72660 123267 72664
rect 123201 72659 123267 72660
rect 124213 72724 124279 72725
rect 124213 72720 124260 72724
rect 124324 72722 124330 72724
rect 124489 72722 124555 72725
rect 124622 72722 124628 72724
rect 124213 72664 124218 72720
rect 124213 72660 124260 72664
rect 124324 72662 124370 72722
rect 124489 72720 124628 72722
rect 124489 72664 124494 72720
rect 124550 72664 124628 72720
rect 124489 72662 124628 72664
rect 124324 72660 124330 72662
rect 124213 72659 124279 72660
rect 124489 72659 124555 72662
rect 124622 72660 124628 72662
rect 124692 72660 124698 72724
rect 125593 72722 125659 72725
rect 125726 72722 125732 72724
rect 125593 72720 125732 72722
rect 125593 72664 125598 72720
rect 125654 72664 125732 72720
rect 125593 72662 125732 72664
rect 125593 72659 125659 72662
rect 125726 72660 125732 72662
rect 125796 72660 125802 72724
rect 25497 72584 103530 72586
rect 25497 72528 25502 72584
rect 25558 72528 103530 72584
rect 25497 72526 103530 72528
rect 117865 72586 117931 72589
rect 123385 72586 123451 72589
rect 123753 72588 123819 72589
rect 117865 72584 123451 72586
rect 117865 72528 117870 72584
rect 117926 72528 123390 72584
rect 123446 72528 123451 72584
rect 117865 72526 123451 72528
rect 25497 72523 25563 72526
rect 117865 72523 117931 72526
rect 123385 72523 123451 72526
rect 123702 72524 123708 72588
rect 123772 72586 123819 72588
rect 124397 72586 124463 72589
rect 124806 72586 124812 72588
rect 123772 72584 123864 72586
rect 123814 72528 123864 72584
rect 123772 72526 123864 72528
rect 124397 72584 124812 72586
rect 124397 72528 124402 72584
rect 124458 72528 124812 72584
rect 124397 72526 124812 72528
rect 123772 72524 123819 72526
rect 123753 72523 123819 72524
rect 124397 72523 124463 72526
rect 124806 72524 124812 72526
rect 124876 72524 124882 72588
rect 126421 72586 126487 72589
rect 126654 72586 126714 72931
rect 126973 72858 127039 72861
rect 127382 72858 127388 72860
rect 126973 72856 127388 72858
rect 126973 72800 126978 72856
rect 127034 72800 127388 72856
rect 126973 72798 127388 72800
rect 126973 72795 127039 72798
rect 127382 72796 127388 72798
rect 127452 72796 127458 72860
rect 128353 72858 128419 72861
rect 128670 72858 128676 72860
rect 128353 72856 128676 72858
rect 128353 72800 128358 72856
rect 128414 72800 128676 72856
rect 128353 72798 128676 72800
rect 128353 72795 128419 72798
rect 128670 72796 128676 72798
rect 128740 72796 128746 72860
rect 129782 72725 129842 73067
rect 130878 72932 130884 72996
rect 130948 72994 130954 72996
rect 134057 72994 134123 72997
rect 130948 72992 134123 72994
rect 130948 72936 134062 72992
rect 134118 72936 134123 72992
rect 130948 72934 134123 72936
rect 130948 72932 130954 72934
rect 134057 72931 134123 72934
rect 142838 72932 142844 72996
rect 142908 72994 142914 72996
rect 143349 72994 143415 72997
rect 142908 72992 143415 72994
rect 142908 72936 143354 72992
rect 143410 72936 143415 72992
rect 142908 72934 143415 72936
rect 142908 72932 142914 72934
rect 143349 72931 143415 72934
rect 145373 72994 145439 72997
rect 145373 72992 147506 72994
rect 145373 72936 145378 72992
rect 145434 72936 147506 72992
rect 145373 72934 147506 72936
rect 145373 72931 145439 72934
rect 131982 72796 131988 72860
rect 132052 72858 132058 72860
rect 132401 72858 132467 72861
rect 132052 72856 132467 72858
rect 132052 72800 132406 72856
rect 132462 72800 132467 72856
rect 132052 72798 132467 72800
rect 132052 72796 132058 72798
rect 132401 72795 132467 72798
rect 133270 72796 133276 72860
rect 133340 72858 133346 72860
rect 133689 72858 133755 72861
rect 133340 72856 133755 72858
rect 133340 72800 133694 72856
rect 133750 72800 133755 72856
rect 133340 72798 133755 72800
rect 133340 72796 133346 72798
rect 133689 72795 133755 72798
rect 135069 72860 135135 72861
rect 135069 72856 135116 72860
rect 135180 72858 135186 72860
rect 136449 72858 136515 72861
rect 136582 72858 136588 72860
rect 135069 72800 135074 72856
rect 135069 72796 135116 72800
rect 135180 72798 135226 72858
rect 136449 72856 136588 72858
rect 136449 72800 136454 72856
rect 136510 72800 136588 72856
rect 136449 72798 136588 72800
rect 135180 72796 135186 72798
rect 135069 72795 135135 72796
rect 136449 72795 136515 72798
rect 136582 72796 136588 72798
rect 136652 72796 136658 72860
rect 137318 72796 137324 72860
rect 137388 72858 137394 72860
rect 137921 72858 137987 72861
rect 137388 72856 137987 72858
rect 137388 72800 137926 72856
rect 137982 72800 137987 72856
rect 137388 72798 137987 72800
rect 137388 72796 137394 72798
rect 137921 72795 137987 72798
rect 143257 72858 143323 72861
rect 143390 72858 143396 72860
rect 143257 72856 143396 72858
rect 143257 72800 143262 72856
rect 143318 72800 143396 72856
rect 143257 72798 143396 72800
rect 143257 72795 143323 72798
rect 143390 72796 143396 72798
rect 143460 72796 143466 72860
rect 144494 72796 144500 72860
rect 144564 72858 144570 72860
rect 144821 72858 144887 72861
rect 144564 72856 144887 72858
rect 144564 72800 144826 72856
rect 144882 72800 144887 72856
rect 144564 72798 144887 72800
rect 144564 72796 144570 72798
rect 144821 72795 144887 72798
rect 145046 72796 145052 72860
rect 145116 72858 145122 72860
rect 146201 72858 146267 72861
rect 145116 72856 146267 72858
rect 145116 72800 146206 72856
rect 146262 72800 146267 72856
rect 145116 72798 146267 72800
rect 147446 72858 147506 72934
rect 147622 72932 147628 72996
rect 147692 72994 147698 72996
rect 147765 72994 147831 72997
rect 153101 72994 153167 72997
rect 147692 72992 147831 72994
rect 147692 72936 147770 72992
rect 147826 72936 147831 72992
rect 147692 72934 147831 72936
rect 147692 72932 147698 72934
rect 147765 72931 147831 72934
rect 148182 72992 153167 72994
rect 148182 72936 153106 72992
rect 153162 72936 153167 72992
rect 148182 72934 153167 72936
rect 148182 72858 148242 72934
rect 153101 72931 153167 72934
rect 153285 72994 153351 72997
rect 153285 72992 156522 72994
rect 153285 72936 153290 72992
rect 153346 72936 156522 72992
rect 153285 72934 156522 72936
rect 153285 72931 153351 72934
rect 147446 72798 148242 72858
rect 145116 72796 145122 72798
rect 146201 72795 146267 72798
rect 148358 72796 148364 72860
rect 148428 72858 148434 72860
rect 148869 72858 148935 72861
rect 148428 72856 148935 72858
rect 148428 72800 148874 72856
rect 148930 72800 148935 72856
rect 148428 72798 148935 72800
rect 148428 72796 148434 72798
rect 148869 72795 148935 72798
rect 150157 72858 150223 72861
rect 150382 72858 150388 72860
rect 150157 72856 150388 72858
rect 150157 72800 150162 72856
rect 150218 72800 150388 72856
rect 150157 72798 150388 72800
rect 150157 72795 150223 72798
rect 150382 72796 150388 72798
rect 150452 72796 150458 72860
rect 152222 72796 152228 72860
rect 152292 72858 152298 72860
rect 152733 72858 152799 72861
rect 152292 72856 152799 72858
rect 152292 72800 152738 72856
rect 152794 72800 152799 72856
rect 152292 72798 152799 72800
rect 152292 72796 152298 72798
rect 152733 72795 152799 72798
rect 153878 72796 153884 72860
rect 153948 72858 153954 72860
rect 154205 72858 154271 72861
rect 153948 72856 154271 72858
rect 153948 72800 154210 72856
rect 154266 72800 154271 72856
rect 153948 72798 154271 72800
rect 153948 72796 153954 72798
rect 154205 72795 154271 72798
rect 155350 72796 155356 72860
rect 155420 72858 155426 72860
rect 155585 72858 155651 72861
rect 155420 72856 155651 72858
rect 155420 72800 155590 72856
rect 155646 72800 155651 72856
rect 155420 72798 155651 72800
rect 155420 72796 155426 72798
rect 155585 72795 155651 72798
rect 127249 72724 127315 72725
rect 127198 72722 127204 72724
rect 127158 72662 127204 72722
rect 127268 72720 127315 72724
rect 127310 72664 127315 72720
rect 127198 72660 127204 72662
rect 127268 72660 127315 72664
rect 128486 72660 128492 72724
rect 128556 72722 128562 72724
rect 128629 72722 128695 72725
rect 128556 72720 128695 72722
rect 128556 72664 128634 72720
rect 128690 72664 128695 72720
rect 128556 72662 128695 72664
rect 129782 72720 129891 72725
rect 129782 72664 129830 72720
rect 129886 72664 129891 72720
rect 129782 72662 129891 72664
rect 128556 72660 128562 72662
rect 127249 72659 127315 72660
rect 128629 72659 128695 72662
rect 129825 72659 129891 72662
rect 132309 72724 132375 72725
rect 133597 72724 133663 72725
rect 134885 72724 134951 72725
rect 136357 72724 136423 72725
rect 132309 72720 132356 72724
rect 132420 72722 132426 72724
rect 132309 72664 132314 72720
rect 132309 72660 132356 72664
rect 132420 72662 132466 72722
rect 133597 72720 133644 72724
rect 133708 72722 133714 72724
rect 133597 72664 133602 72720
rect 132420 72660 132426 72662
rect 133597 72660 133644 72664
rect 133708 72662 133754 72722
rect 134885 72720 134932 72724
rect 134996 72722 135002 72724
rect 134885 72664 134890 72720
rect 133708 72660 133714 72662
rect 134885 72660 134932 72664
rect 134996 72662 135042 72722
rect 136357 72720 136404 72724
rect 136468 72722 136474 72724
rect 136357 72664 136362 72720
rect 134996 72660 135002 72662
rect 136357 72660 136404 72664
rect 136468 72662 136514 72722
rect 136468 72660 136474 72662
rect 137502 72660 137508 72724
rect 137572 72722 137578 72724
rect 137829 72722 137895 72725
rect 137572 72720 137895 72722
rect 137572 72664 137834 72720
rect 137890 72664 137895 72720
rect 137572 72662 137895 72664
rect 137572 72660 137578 72662
rect 132309 72659 132375 72660
rect 133597 72659 133663 72660
rect 134885 72659 134951 72660
rect 136357 72659 136423 72660
rect 137829 72659 137895 72662
rect 143022 72660 143028 72724
rect 143092 72722 143098 72724
rect 143165 72722 143231 72725
rect 143092 72720 143231 72722
rect 143092 72664 143170 72720
rect 143226 72664 143231 72720
rect 143092 72662 143231 72664
rect 143092 72660 143098 72662
rect 143165 72659 143231 72662
rect 144729 72722 144795 72725
rect 146109 72724 146175 72725
rect 144862 72722 144868 72724
rect 144729 72720 144868 72722
rect 144729 72664 144734 72720
rect 144790 72664 144868 72720
rect 144729 72662 144868 72664
rect 144729 72659 144795 72662
rect 144862 72660 144868 72662
rect 144932 72660 144938 72724
rect 146109 72720 146156 72724
rect 146220 72722 146226 72724
rect 146109 72664 146114 72720
rect 146109 72660 146156 72664
rect 146220 72662 146266 72722
rect 146220 72660 146226 72662
rect 147070 72660 147076 72724
rect 147140 72722 147146 72724
rect 147305 72722 147371 72725
rect 147140 72720 147371 72722
rect 147140 72664 147310 72720
rect 147366 72664 147371 72720
rect 147140 72662 147371 72664
rect 147140 72660 147146 72662
rect 146109 72659 146175 72660
rect 147305 72659 147371 72662
rect 147630 72662 148058 72722
rect 126421 72584 126714 72586
rect 126421 72528 126426 72584
rect 126482 72528 126714 72584
rect 126421 72526 126714 72528
rect 127157 72586 127223 72589
rect 127566 72586 127572 72588
rect 127157 72584 127572 72586
rect 127157 72528 127162 72584
rect 127218 72528 127572 72584
rect 127157 72526 127572 72528
rect 126421 72523 126487 72526
rect 127157 72523 127223 72526
rect 127566 72524 127572 72526
rect 127636 72524 127642 72588
rect 128445 72586 128511 72589
rect 128854 72586 128860 72588
rect 128445 72584 128860 72586
rect 128445 72528 128450 72584
rect 128506 72528 128860 72584
rect 128445 72526 128860 72528
rect 128445 72523 128511 72526
rect 128854 72524 128860 72526
rect 128924 72524 128930 72588
rect 133086 72524 133092 72588
rect 133156 72586 133162 72588
rect 133505 72586 133571 72589
rect 133156 72584 133571 72586
rect 133156 72528 133510 72584
rect 133566 72528 133571 72584
rect 133156 72526 133571 72528
rect 133156 72524 133162 72526
rect 133505 72523 133571 72526
rect 134742 72524 134748 72588
rect 134812 72586 134818 72588
rect 135161 72586 135227 72589
rect 134812 72584 135227 72586
rect 134812 72528 135166 72584
rect 135222 72528 135227 72584
rect 134812 72526 135227 72528
rect 134812 72524 134818 72526
rect 135161 72523 135227 72526
rect 136214 72524 136220 72588
rect 136284 72586 136290 72588
rect 136541 72586 136607 72589
rect 136284 72584 136607 72586
rect 136284 72528 136546 72584
rect 136602 72528 136607 72584
rect 136284 72526 136607 72528
rect 136284 72524 136290 72526
rect 136541 72523 136607 72526
rect 143206 72524 143212 72588
rect 143276 72586 143282 72588
rect 143441 72586 143507 72589
rect 143276 72584 143507 72586
rect 143276 72528 143446 72584
rect 143502 72528 143507 72584
rect 143276 72526 143507 72528
rect 143276 72524 143282 72526
rect 143441 72523 143507 72526
rect 144310 72524 144316 72588
rect 144380 72586 144386 72588
rect 144637 72586 144703 72589
rect 144380 72584 144703 72586
rect 144380 72528 144642 72584
rect 144698 72528 144703 72584
rect 144380 72526 144703 72528
rect 144380 72524 144386 72526
rect 144637 72523 144703 72526
rect 144821 72586 144887 72589
rect 147630 72586 147690 72662
rect 144821 72584 147690 72586
rect 144821 72528 144826 72584
rect 144882 72528 147690 72584
rect 144821 72526 147690 72528
rect 144821 72523 144887 72526
rect 122833 72450 122899 72453
rect 123334 72450 123340 72452
rect 122833 72448 123340 72450
rect 122833 72392 122838 72448
rect 122894 72392 123340 72448
rect 122833 72390 123340 72392
rect 122833 72387 122899 72390
rect 123334 72388 123340 72390
rect 123404 72388 123410 72452
rect 127014 72388 127020 72452
rect 127084 72450 127090 72452
rect 127341 72450 127407 72453
rect 127084 72448 127407 72450
rect 127084 72392 127346 72448
rect 127402 72392 127407 72448
rect 127084 72390 127407 72392
rect 127084 72388 127090 72390
rect 127341 72387 127407 72390
rect 133454 72388 133460 72452
rect 133524 72450 133530 72452
rect 133781 72450 133847 72453
rect 133524 72448 133847 72450
rect 133524 72392 133786 72448
rect 133842 72392 133847 72448
rect 133524 72390 133847 72392
rect 133524 72388 133530 72390
rect 133781 72387 133847 72390
rect 134558 72388 134564 72452
rect 134628 72450 134634 72452
rect 134793 72450 134859 72453
rect 134628 72448 134859 72450
rect 134628 72392 134798 72448
rect 134854 72392 134859 72448
rect 134628 72390 134859 72392
rect 134628 72388 134634 72390
rect 134793 72387 134859 72390
rect 136030 72388 136036 72452
rect 136100 72450 136106 72452
rect 136265 72450 136331 72453
rect 139577 72450 139643 72453
rect 136100 72448 136331 72450
rect 136100 72392 136270 72448
rect 136326 72392 136331 72448
rect 136100 72390 136331 72392
rect 136100 72388 136106 72390
rect 136265 72387 136331 72390
rect 136406 72448 139643 72450
rect 136406 72392 139582 72448
rect 139638 72392 139643 72448
rect 136406 72390 139643 72392
rect 132166 72252 132172 72316
rect 132236 72314 132242 72316
rect 136406 72314 136466 72390
rect 139577 72387 139643 72390
rect 144126 72388 144132 72452
rect 144196 72450 144202 72452
rect 144545 72450 144611 72453
rect 144196 72448 144611 72450
rect 144196 72392 144550 72448
rect 144606 72392 144611 72448
rect 144196 72390 144611 72392
rect 147998 72450 148058 72662
rect 148542 72660 148548 72724
rect 148612 72722 148618 72724
rect 148777 72722 148843 72725
rect 148612 72720 148843 72722
rect 148612 72664 148782 72720
rect 148838 72664 148843 72720
rect 148612 72662 148843 72664
rect 148612 72660 148618 72662
rect 148777 72659 148843 72662
rect 150198 72660 150204 72724
rect 150268 72722 150274 72724
rect 150341 72722 150407 72725
rect 150268 72720 150407 72722
rect 150268 72664 150346 72720
rect 150402 72664 150407 72720
rect 150268 72662 150407 72664
rect 150268 72660 150274 72662
rect 150341 72659 150407 72662
rect 151537 72722 151603 72725
rect 151670 72722 151676 72724
rect 151537 72720 151676 72722
rect 151537 72664 151542 72720
rect 151598 72664 151676 72720
rect 151537 72662 151676 72664
rect 151537 72659 151603 72662
rect 151670 72660 151676 72662
rect 151740 72660 151746 72724
rect 152406 72660 152412 72724
rect 152476 72722 152482 72724
rect 153009 72722 153075 72725
rect 154297 72724 154363 72725
rect 155769 72724 155835 72725
rect 154246 72722 154252 72724
rect 152476 72720 153075 72722
rect 152476 72664 153014 72720
rect 153070 72664 153075 72720
rect 152476 72662 153075 72664
rect 154206 72662 154252 72722
rect 154316 72720 154363 72724
rect 155718 72722 155724 72724
rect 154358 72664 154363 72720
rect 152476 72660 152482 72662
rect 153009 72659 153075 72662
rect 154246 72660 154252 72662
rect 154316 72660 154363 72664
rect 155678 72662 155724 72722
rect 155788 72720 155835 72724
rect 155830 72664 155835 72720
rect 155718 72660 155724 72662
rect 155788 72660 155835 72664
rect 156462 72722 156522 72934
rect 157382 72858 157442 73070
rect 157517 73128 157564 73132
rect 157628 73130 157634 73132
rect 157977 73130 158043 73133
rect 161430 73130 161490 73206
rect 157517 73072 157522 73128
rect 157517 73068 157564 73072
rect 157628 73070 157674 73130
rect 157977 73128 161490 73130
rect 157977 73072 157982 73128
rect 158038 73072 161490 73128
rect 157977 73070 161490 73072
rect 157628 73068 157634 73070
rect 157517 73067 157583 73068
rect 157977 73067 158043 73070
rect 162158 73068 162164 73132
rect 162228 73130 162234 73132
rect 162577 73130 162643 73133
rect 162228 73128 162643 73130
rect 162228 73072 162582 73128
rect 162638 73072 162643 73128
rect 162228 73070 162643 73072
rect 164190 73130 164250 73206
rect 169109 73130 169175 73133
rect 164190 73128 169175 73130
rect 164190 73072 169114 73128
rect 169170 73072 169175 73128
rect 164190 73070 169175 73072
rect 162228 73068 162234 73070
rect 162577 73067 162643 73070
rect 169109 73067 169175 73070
rect 159030 72932 159036 72996
rect 159100 72994 159106 72996
rect 169109 72994 169175 72997
rect 159100 72992 169175 72994
rect 159100 72936 169114 72992
rect 169170 72936 169175 72992
rect 159100 72934 169175 72936
rect 159100 72932 159106 72934
rect 169109 72931 169175 72934
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 169201 72858 169267 72861
rect 157382 72856 169267 72858
rect 157382 72800 169206 72856
rect 169262 72800 169267 72856
rect 583520 72844 584960 72934
rect 157382 72798 169267 72800
rect 169201 72795 169267 72798
rect 157977 72722 158043 72725
rect 158345 72724 158411 72725
rect 158294 72722 158300 72724
rect 156462 72720 158043 72722
rect 156462 72664 157982 72720
rect 158038 72664 158043 72720
rect 156462 72662 158043 72664
rect 158254 72662 158300 72722
rect 158364 72720 158411 72724
rect 158406 72664 158411 72720
rect 154297 72659 154363 72660
rect 155769 72659 155835 72660
rect 157977 72659 158043 72662
rect 158294 72660 158300 72662
rect 158364 72660 158411 72664
rect 158345 72659 158411 72660
rect 158529 72722 158595 72725
rect 159173 72724 159239 72725
rect 159633 72724 159699 72725
rect 158662 72722 158668 72724
rect 158529 72720 158668 72722
rect 158529 72664 158534 72720
rect 158590 72664 158668 72720
rect 158529 72662 158668 72664
rect 158529 72659 158595 72662
rect 158662 72660 158668 72662
rect 158732 72660 158738 72724
rect 159173 72720 159220 72724
rect 159284 72722 159290 72724
rect 159582 72722 159588 72724
rect 159173 72664 159178 72720
rect 159173 72660 159220 72664
rect 159284 72662 159330 72722
rect 159542 72662 159588 72722
rect 159652 72720 159699 72724
rect 159694 72664 159699 72720
rect 159284 72660 159290 72662
rect 159582 72660 159588 72662
rect 159652 72660 159699 72664
rect 159766 72660 159772 72724
rect 159836 72722 159842 72724
rect 159909 72722 159975 72725
rect 159836 72720 159975 72722
rect 159836 72664 159914 72720
rect 159970 72664 159975 72720
rect 159836 72662 159975 72664
rect 159836 72660 159842 72662
rect 159173 72659 159239 72660
rect 159633 72659 159699 72660
rect 159909 72659 159975 72662
rect 160277 72722 160343 72725
rect 161013 72722 161079 72725
rect 160277 72720 161079 72722
rect 160277 72664 160282 72720
rect 160338 72664 161018 72720
rect 161074 72664 161079 72720
rect 160277 72662 161079 72664
rect 160277 72659 160343 72662
rect 161013 72659 161079 72662
rect 162526 72660 162532 72724
rect 162596 72722 162602 72724
rect 162669 72722 162735 72725
rect 162596 72720 162735 72722
rect 162596 72664 162674 72720
rect 162730 72664 162735 72720
rect 162596 72662 162735 72664
rect 162596 72660 162602 72662
rect 162669 72659 162735 72662
rect 163446 72660 163452 72724
rect 163516 72722 163522 72724
rect 164141 72722 164207 72725
rect 165337 72724 165403 72725
rect 165286 72722 165292 72724
rect 163516 72720 164207 72722
rect 163516 72664 164146 72720
rect 164202 72664 164207 72720
rect 163516 72662 164207 72664
rect 165246 72662 165292 72722
rect 165356 72720 165403 72724
rect 332593 72722 332659 72725
rect 165398 72664 165403 72720
rect 163516 72660 163522 72662
rect 164141 72659 164207 72662
rect 165286 72660 165292 72662
rect 165356 72660 165403 72664
rect 165337 72659 165403 72660
rect 166398 72720 332659 72722
rect 166398 72664 332598 72720
rect 332654 72664 332659 72720
rect 166398 72662 332659 72664
rect 148174 72524 148180 72588
rect 148244 72586 148250 72588
rect 148961 72586 149027 72589
rect 148244 72584 149027 72586
rect 148244 72528 148966 72584
rect 149022 72528 149027 72584
rect 148244 72526 149027 72528
rect 148244 72524 148250 72526
rect 148961 72523 149027 72526
rect 151118 72524 151124 72588
rect 151188 72586 151194 72588
rect 151445 72586 151511 72589
rect 151188 72584 151511 72586
rect 151188 72528 151450 72584
rect 151506 72528 151511 72584
rect 151188 72526 151511 72528
rect 151188 72524 151194 72526
rect 151445 72523 151511 72526
rect 154062 72524 154068 72588
rect 154132 72586 154138 72588
rect 154481 72586 154547 72589
rect 154132 72584 154547 72586
rect 154132 72528 154486 72584
rect 154542 72528 154547 72584
rect 154132 72526 154547 72528
rect 154132 72524 154138 72526
rect 154481 72523 154547 72526
rect 155166 72524 155172 72588
rect 155236 72586 155242 72588
rect 155677 72586 155743 72589
rect 157241 72588 157307 72589
rect 157190 72586 157196 72588
rect 155236 72584 155743 72586
rect 155236 72528 155682 72584
rect 155738 72528 155743 72584
rect 155236 72526 155743 72528
rect 157150 72526 157196 72586
rect 157260 72584 157307 72588
rect 157302 72528 157307 72584
rect 155236 72524 155242 72526
rect 155677 72523 155743 72526
rect 157190 72524 157196 72526
rect 157260 72524 157307 72528
rect 157926 72524 157932 72588
rect 157996 72586 158002 72588
rect 158621 72586 158687 72589
rect 157996 72584 158687 72586
rect 157996 72528 158626 72584
rect 158682 72528 158687 72584
rect 157996 72526 158687 72528
rect 157996 72524 158002 72526
rect 157241 72523 157307 72524
rect 158621 72523 158687 72526
rect 159398 72524 159404 72588
rect 159468 72586 159474 72588
rect 159817 72586 159883 72589
rect 159468 72584 159883 72586
rect 159468 72528 159822 72584
rect 159878 72528 159883 72584
rect 159468 72526 159883 72528
rect 159468 72524 159474 72526
rect 159817 72523 159883 72526
rect 161054 72524 161060 72588
rect 161124 72586 161130 72588
rect 161381 72586 161447 72589
rect 161124 72584 161447 72586
rect 161124 72528 161386 72584
rect 161442 72528 161447 72584
rect 161124 72526 161447 72528
rect 161124 72524 161130 72526
rect 161381 72523 161447 72526
rect 162485 72586 162551 72589
rect 162710 72586 162716 72588
rect 162485 72584 162716 72586
rect 162485 72528 162490 72584
rect 162546 72528 162716 72584
rect 162485 72526 162716 72528
rect 162485 72523 162551 72526
rect 162710 72524 162716 72526
rect 162780 72524 162786 72588
rect 163957 72586 164023 72589
rect 164141 72586 164207 72589
rect 163957 72584 164207 72586
rect 163957 72528 163962 72584
rect 164018 72528 164146 72584
rect 164202 72528 164207 72584
rect 163957 72526 164207 72528
rect 163957 72523 164023 72526
rect 164141 72523 164207 72526
rect 165429 72588 165495 72589
rect 165429 72584 165476 72588
rect 165540 72586 165546 72588
rect 165705 72586 165771 72589
rect 166398 72586 166458 72662
rect 332593 72659 332659 72662
rect 165429 72528 165434 72584
rect 165429 72524 165476 72528
rect 165540 72526 165586 72586
rect 165705 72584 166458 72586
rect 165705 72528 165710 72584
rect 165766 72528 166458 72584
rect 165705 72526 166458 72528
rect 166533 72588 166599 72589
rect 166533 72584 166580 72588
rect 166644 72586 166650 72588
rect 501781 72586 501847 72589
rect 166533 72528 166538 72584
rect 165540 72524 165546 72526
rect 165429 72523 165495 72524
rect 165705 72523 165771 72526
rect 166533 72524 166580 72528
rect 166644 72526 166690 72586
rect 166950 72584 501847 72586
rect 166950 72528 501786 72584
rect 501842 72528 501847 72584
rect 166950 72526 501847 72528
rect 166644 72524 166650 72526
rect 166533 72523 166599 72524
rect 151077 72450 151143 72453
rect 147998 72448 151143 72450
rect 147998 72392 151082 72448
rect 151138 72392 151143 72448
rect 147998 72390 151143 72392
rect 144196 72388 144202 72390
rect 144545 72387 144611 72390
rect 151077 72387 151143 72390
rect 151302 72388 151308 72452
rect 151372 72450 151378 72452
rect 151721 72450 151787 72453
rect 151372 72448 151787 72450
rect 151372 72392 151726 72448
rect 151782 72392 151787 72448
rect 151372 72390 151787 72392
rect 151372 72388 151378 72390
rect 151721 72387 151787 72390
rect 154113 72450 154179 72453
rect 154430 72450 154436 72452
rect 154113 72448 154436 72450
rect 154113 72392 154118 72448
rect 154174 72392 154436 72448
rect 154113 72390 154436 72392
rect 154113 72387 154179 72390
rect 154430 72388 154436 72390
rect 154500 72388 154506 72452
rect 155534 72388 155540 72452
rect 155604 72450 155610 72452
rect 155861 72450 155927 72453
rect 155604 72448 155927 72450
rect 155604 72392 155866 72448
rect 155922 72392 155927 72448
rect 155604 72390 155927 72392
rect 155604 72388 155610 72390
rect 155861 72387 155927 72390
rect 156646 72390 157350 72450
rect 132236 72254 136466 72314
rect 136817 72314 136883 72317
rect 142061 72314 142127 72317
rect 143717 72314 143783 72317
rect 136817 72312 138030 72314
rect 136817 72256 136822 72312
rect 136878 72256 138030 72312
rect 136817 72254 138030 72256
rect 132236 72252 132242 72254
rect 136817 72251 136883 72254
rect 116853 72042 116919 72045
rect 122373 72042 122439 72045
rect 116853 72040 122439 72042
rect 116853 71984 116858 72040
rect 116914 71984 122378 72040
rect 122434 71984 122439 72040
rect 116853 71982 122439 71984
rect 137970 72042 138030 72254
rect 142061 72312 143783 72314
rect 142061 72256 142066 72312
rect 142122 72256 143722 72312
rect 143778 72256 143783 72312
rect 142061 72254 143783 72256
rect 142061 72251 142127 72254
rect 143717 72251 143783 72254
rect 153837 72314 153903 72317
rect 156137 72314 156203 72317
rect 153837 72312 156203 72314
rect 153837 72256 153842 72312
rect 153898 72256 156142 72312
rect 156198 72256 156203 72312
rect 153837 72254 156203 72256
rect 153837 72251 153903 72254
rect 156137 72251 156203 72254
rect 138473 72178 138539 72181
rect 144821 72178 144887 72181
rect 138473 72176 144887 72178
rect 138473 72120 138478 72176
rect 138534 72120 144826 72176
rect 144882 72120 144887 72176
rect 138473 72118 144887 72120
rect 138473 72115 138539 72118
rect 144821 72115 144887 72118
rect 146886 72116 146892 72180
rect 146956 72178 146962 72180
rect 147397 72178 147463 72181
rect 146956 72176 147463 72178
rect 146956 72120 147402 72176
rect 147458 72120 147463 72176
rect 146956 72118 147463 72120
rect 146956 72116 146962 72118
rect 147397 72115 147463 72118
rect 147765 72178 147831 72181
rect 156646 72178 156706 72390
rect 157290 72314 157350 72390
rect 157742 72388 157748 72452
rect 157812 72450 157818 72452
rect 158437 72450 158503 72453
rect 157812 72448 158503 72450
rect 157812 72392 158442 72448
rect 158498 72392 158503 72448
rect 157812 72390 158503 72392
rect 157812 72388 157818 72390
rect 158437 72387 158503 72390
rect 158621 72450 158687 72453
rect 159030 72450 159036 72452
rect 158621 72448 159036 72450
rect 158621 72392 158626 72448
rect 158682 72392 159036 72448
rect 158621 72390 159036 72392
rect 158621 72387 158687 72390
rect 159030 72388 159036 72390
rect 159100 72388 159106 72452
rect 160553 72450 160619 72453
rect 160553 72448 162226 72450
rect 160553 72392 160558 72448
rect 160614 72392 162226 72448
rect 160553 72390 162226 72392
rect 160553 72387 160619 72390
rect 161422 72314 161428 72316
rect 157290 72254 161428 72314
rect 161422 72252 161428 72254
rect 161492 72252 161498 72316
rect 162166 72314 162226 72390
rect 162342 72388 162348 72452
rect 162412 72450 162418 72452
rect 162761 72450 162827 72453
rect 162412 72448 162827 72450
rect 162412 72392 162766 72448
rect 162822 72392 162827 72448
rect 162412 72390 162827 72392
rect 162412 72388 162418 72390
rect 162761 72387 162827 72390
rect 163078 72388 163084 72452
rect 163148 72450 163154 72452
rect 164049 72450 164115 72453
rect 163148 72448 164115 72450
rect 163148 72392 164054 72448
rect 164110 72392 164115 72448
rect 163148 72390 164115 72392
rect 163148 72388 163154 72390
rect 164049 72387 164115 72390
rect 165102 72388 165108 72452
rect 165172 72450 165178 72452
rect 165521 72450 165587 72453
rect 165172 72448 165587 72450
rect 165172 72392 165526 72448
rect 165582 72392 165587 72448
rect 165172 72390 165587 72392
rect 165172 72388 165178 72390
rect 165521 72387 165587 72390
rect 166441 72450 166507 72453
rect 166758 72450 166764 72452
rect 166441 72448 166764 72450
rect 166441 72392 166446 72448
rect 166502 72392 166764 72448
rect 166441 72390 166764 72392
rect 166441 72387 166507 72390
rect 166758 72388 166764 72390
rect 166828 72388 166834 72452
rect 166950 72314 167010 72526
rect 501781 72523 501847 72526
rect 162166 72254 167010 72314
rect 168281 72314 168347 72317
rect 178953 72314 179019 72317
rect 168281 72312 179019 72314
rect 168281 72256 168286 72312
rect 168342 72256 178958 72312
rect 179014 72256 179019 72312
rect 168281 72254 179019 72256
rect 168281 72251 168347 72254
rect 178953 72251 179019 72254
rect 147765 72176 156706 72178
rect 147765 72120 147770 72176
rect 147826 72120 156706 72176
rect 147765 72118 156706 72120
rect 147765 72115 147831 72118
rect 157558 72116 157564 72180
rect 157628 72178 157634 72180
rect 157977 72178 158043 72181
rect 157628 72176 158043 72178
rect 157628 72120 157982 72176
rect 158038 72120 158043 72176
rect 157628 72118 158043 72120
rect 157628 72116 157634 72118
rect 157977 72115 158043 72118
rect 158345 72178 158411 72181
rect 165705 72178 165771 72181
rect 158345 72176 165771 72178
rect 158345 72120 158350 72176
rect 158406 72120 165710 72176
rect 165766 72120 165771 72176
rect 158345 72118 165771 72120
rect 158345 72115 158411 72118
rect 165705 72115 165771 72118
rect 166349 72180 166415 72181
rect 166349 72176 166396 72180
rect 166460 72178 166466 72180
rect 166625 72178 166691 72181
rect 167494 72178 167500 72180
rect 166349 72120 166354 72176
rect 166349 72116 166396 72120
rect 166460 72118 166506 72178
rect 166625 72176 167500 72178
rect 166625 72120 166630 72176
rect 166686 72120 167500 72176
rect 166625 72118 167500 72120
rect 166460 72116 166466 72118
rect 166349 72115 166415 72116
rect 166625 72115 166691 72118
rect 167494 72116 167500 72118
rect 167564 72116 167570 72180
rect 160870 72042 160876 72044
rect 137970 71982 160876 72042
rect 116853 71979 116919 71982
rect 122373 71979 122439 71982
rect 160870 71980 160876 71982
rect 160940 71980 160946 72044
rect 166717 72042 166783 72045
rect 166717 72040 176670 72042
rect 166717 71984 166722 72040
rect 166778 71984 176670 72040
rect 166717 71982 176670 71984
rect 166717 71979 166783 71982
rect 138197 71906 138263 71909
rect 147622 71906 147628 71908
rect 138197 71904 147628 71906
rect 138197 71848 138202 71904
rect 138258 71848 147628 71904
rect 138197 71846 147628 71848
rect 138197 71843 138263 71846
rect 147622 71844 147628 71846
rect 147692 71844 147698 71908
rect 151077 71906 151143 71909
rect 155902 71906 155908 71908
rect 151077 71904 155908 71906
rect 151077 71848 151082 71904
rect 151138 71848 155908 71904
rect 151077 71846 155908 71848
rect 151077 71843 151143 71846
rect 155902 71844 155908 71846
rect 155972 71844 155978 71908
rect 156086 71844 156092 71908
rect 156156 71906 156162 71908
rect 157149 71906 157215 71909
rect 156156 71904 157215 71906
rect 156156 71848 157154 71904
rect 157210 71848 157215 71904
rect 156156 71846 157215 71848
rect 156156 71844 156162 71846
rect 157149 71843 157215 71846
rect 163313 71906 163379 71909
rect 165705 71906 165771 71909
rect 163313 71904 165771 71906
rect 163313 71848 163318 71904
rect 163374 71848 165710 71904
rect 165766 71848 165771 71904
rect 163313 71846 165771 71848
rect 163313 71843 163379 71846
rect 165705 71843 165771 71846
rect 166206 71844 166212 71908
rect 166276 71906 166282 71908
rect 170489 71906 170555 71909
rect 166276 71904 170555 71906
rect 166276 71848 170494 71904
rect 170550 71848 170555 71904
rect 166276 71846 170555 71848
rect 176610 71906 176670 71982
rect 577497 71906 577563 71909
rect 176610 71904 577563 71906
rect 176610 71848 577502 71904
rect 577558 71848 577563 71904
rect 176610 71846 577563 71848
rect 166276 71844 166282 71846
rect 170489 71843 170555 71846
rect 577497 71843 577563 71846
rect 120073 71770 120139 71773
rect 168373 71770 168439 71773
rect 120073 71768 168439 71770
rect -960 71634 480 71724
rect 120073 71712 120078 71768
rect 120134 71712 168378 71768
rect 168434 71712 168439 71768
rect 120073 71710 168439 71712
rect 120073 71707 120139 71710
rect 168373 71707 168439 71710
rect 168281 71634 168347 71637
rect 580349 71634 580415 71637
rect -960 71632 168347 71634
rect -960 71576 168286 71632
rect 168342 71576 168347 71632
rect -960 71574 168347 71576
rect -960 71484 480 71574
rect 168281 71571 168347 71574
rect 171918 71632 580415 71634
rect 171918 71576 580354 71632
rect 580410 71576 580415 71632
rect 171918 71574 580415 71576
rect 137737 71498 137803 71501
rect 147489 71500 147555 71501
rect 147438 71498 147444 71500
rect 137737 71496 138030 71498
rect 137737 71440 137742 71496
rect 137798 71440 138030 71496
rect 137737 71438 138030 71440
rect 147398 71438 147444 71498
rect 147508 71496 147555 71500
rect 147550 71440 147555 71496
rect 137737 71435 137803 71438
rect 105721 71226 105787 71229
rect 129825 71226 129891 71229
rect 105721 71224 129891 71226
rect 105721 71168 105726 71224
rect 105782 71168 129830 71224
rect 129886 71168 129891 71224
rect 105721 71166 129891 71168
rect 137970 71226 138030 71438
rect 147438 71436 147444 71438
rect 147508 71436 147555 71440
rect 147489 71435 147555 71436
rect 167269 71498 167335 71501
rect 171918 71498 171978 71574
rect 580349 71571 580415 71574
rect 580533 71498 580599 71501
rect 167269 71496 171978 71498
rect 167269 71440 167274 71496
rect 167330 71440 171978 71496
rect 167269 71438 171978 71440
rect 176610 71496 580599 71498
rect 176610 71440 580538 71496
rect 580594 71440 580599 71496
rect 176610 71438 580599 71440
rect 167269 71435 167335 71438
rect 147254 71300 147260 71364
rect 147324 71362 147330 71364
rect 147581 71362 147647 71365
rect 147324 71360 147647 71362
rect 147324 71304 147586 71360
rect 147642 71304 147647 71360
rect 147324 71302 147647 71304
rect 147324 71300 147330 71302
rect 147581 71299 147647 71302
rect 160737 71362 160803 71365
rect 161606 71362 161612 71364
rect 160737 71360 161612 71362
rect 160737 71304 160742 71360
rect 160798 71304 161612 71360
rect 160737 71302 161612 71304
rect 160737 71299 160803 71302
rect 161606 71300 161612 71302
rect 161676 71300 161682 71364
rect 167177 71362 167243 71365
rect 176610 71362 176670 71438
rect 580533 71435 580599 71438
rect 167177 71360 176670 71362
rect 167177 71304 167182 71360
rect 167238 71304 176670 71360
rect 167177 71302 176670 71304
rect 167177 71299 167243 71302
rect 208577 71226 208643 71229
rect 137970 71224 208643 71226
rect 137970 71168 208582 71224
rect 208638 71168 208643 71224
rect 137970 71166 208643 71168
rect 105721 71163 105787 71166
rect 129825 71163 129891 71166
rect 208577 71163 208643 71166
rect 18229 71090 18295 71093
rect 123661 71090 123727 71093
rect 18229 71088 123727 71090
rect 18229 71032 18234 71088
rect 18290 71032 123666 71088
rect 123722 71032 123727 71088
rect 18229 71030 123727 71032
rect 18229 71027 18295 71030
rect 123661 71027 123727 71030
rect 165061 71090 165127 71093
rect 559741 71090 559807 71093
rect 165061 71088 559807 71090
rect 165061 71032 165066 71088
rect 165122 71032 559746 71088
rect 559802 71032 559807 71088
rect 165061 71030 559807 71032
rect 165061 71027 165127 71030
rect 559741 71027 559807 71030
rect 121453 70546 121519 70549
rect 118650 70544 121519 70546
rect 118650 70488 121458 70544
rect 121514 70488 121519 70544
rect 118650 70486 121519 70488
rect 117957 70410 118023 70413
rect 118650 70410 118710 70486
rect 121453 70483 121519 70486
rect 117957 70408 118710 70410
rect 117957 70352 117962 70408
rect 118018 70352 118710 70408
rect 117957 70350 118710 70352
rect 162209 70410 162275 70413
rect 162761 70410 162827 70413
rect 162209 70408 162827 70410
rect 162209 70352 162214 70408
rect 162270 70352 162766 70408
rect 162822 70352 162827 70408
rect 162209 70350 162827 70352
rect 117957 70347 118023 70350
rect 162209 70347 162275 70350
rect 162761 70347 162827 70350
rect 44817 70274 44883 70277
rect 168741 70274 168807 70277
rect 44817 70272 168807 70274
rect 44817 70216 44822 70272
rect 44878 70216 168746 70272
rect 168802 70216 168807 70272
rect 44817 70214 168807 70216
rect 44817 70211 44883 70214
rect 168741 70211 168807 70214
rect 104157 70138 104223 70141
rect 168649 70138 168715 70141
rect 104157 70136 168715 70138
rect 104157 70080 104162 70136
rect 104218 70080 168654 70136
rect 168710 70080 168715 70136
rect 104157 70078 168715 70080
rect 104157 70075 104223 70078
rect 168649 70075 168715 70078
rect 90357 69730 90423 69733
rect 128537 69730 128603 69733
rect 90357 69728 128603 69730
rect 90357 69672 90362 69728
rect 90418 69672 128542 69728
rect 128598 69672 128603 69728
rect 90357 69670 128603 69672
rect 90357 69667 90423 69670
rect 128537 69667 128603 69670
rect 141969 69730 142035 69733
rect 262949 69730 263015 69733
rect 141969 69728 263015 69730
rect 141969 69672 141974 69728
rect 142030 69672 262954 69728
rect 263010 69672 263015 69728
rect 141969 69670 263015 69672
rect 141969 69667 142035 69670
rect 262949 69667 263015 69670
rect 116669 69594 116735 69597
rect 121494 69594 121500 69596
rect 116669 69592 121500 69594
rect 116669 69536 116674 69592
rect 116730 69536 121500 69592
rect 116669 69534 121500 69536
rect 116669 69531 116735 69534
rect 121494 69532 121500 69534
rect 121564 69532 121570 69596
rect 150382 69532 150388 69596
rect 150452 69594 150458 69596
rect 368197 69594 368263 69597
rect 150452 69592 368263 69594
rect 150452 69536 368202 69592
rect 368258 69536 368263 69592
rect 150452 69534 368263 69536
rect 150452 69532 150458 69534
rect 368197 69531 368263 69534
rect 134558 68580 134564 68644
rect 134628 68642 134634 68644
rect 170765 68642 170831 68645
rect 134628 68640 170831 68642
rect 134628 68584 170770 68640
rect 170826 68584 170831 68640
rect 134628 68582 170831 68584
rect 134628 68580 134634 68582
rect 170765 68579 170831 68582
rect 136582 68444 136588 68508
rect 136652 68506 136658 68508
rect 192017 68506 192083 68509
rect 136652 68504 192083 68506
rect 136652 68448 192022 68504
rect 192078 68448 192083 68504
rect 136652 68446 192083 68448
rect 136652 68444 136658 68446
rect 192017 68443 192083 68446
rect 139342 68308 139348 68372
rect 139412 68370 139418 68372
rect 227529 68370 227595 68373
rect 139412 68368 227595 68370
rect 139412 68312 227534 68368
rect 227590 68312 227595 68368
rect 139412 68310 227595 68312
rect 139412 68308 139418 68310
rect 227529 68307 227595 68310
rect 72601 68234 72667 68237
rect 127566 68234 127572 68236
rect 72601 68232 127572 68234
rect 72601 68176 72606 68232
rect 72662 68176 127572 68232
rect 72601 68174 127572 68176
rect 72601 68171 72667 68174
rect 127566 68172 127572 68174
rect 127636 68172 127642 68236
rect 163078 68172 163084 68236
rect 163148 68234 163154 68236
rect 475377 68234 475443 68237
rect 163148 68232 475443 68234
rect 163148 68176 475382 68232
rect 475438 68176 475443 68232
rect 163148 68174 475443 68176
rect 163148 68172 163154 68174
rect 475377 68171 475443 68174
rect 158662 67084 158668 67148
rect 158732 67146 158738 67148
rect 173249 67146 173315 67149
rect 158732 67144 173315 67146
rect 158732 67088 173254 67144
rect 173310 67088 173315 67144
rect 158732 67086 173315 67088
rect 158732 67084 158738 67086
rect 173249 67083 173315 67086
rect 34789 67010 34855 67013
rect 124254 67010 124260 67012
rect 34789 67008 124260 67010
rect 34789 66952 34794 67008
rect 34850 66952 124260 67008
rect 34789 66950 124260 66952
rect 34789 66947 34855 66950
rect 124254 66948 124260 66950
rect 124324 66948 124330 67012
rect 144862 66948 144868 67012
rect 144932 67010 144938 67012
rect 298461 67010 298527 67013
rect 144932 67008 298527 67010
rect 144932 66952 298466 67008
rect 298522 66952 298527 67008
rect 144932 66950 298527 66952
rect 144932 66948 144938 66950
rect 298461 66947 298527 66950
rect 21817 66874 21883 66877
rect 123150 66874 123156 66876
rect 21817 66872 123156 66874
rect 21817 66816 21822 66872
rect 21878 66816 123156 66872
rect 21817 66814 123156 66816
rect 21817 66811 21883 66814
rect 123150 66812 123156 66814
rect 123220 66812 123226 66876
rect 147806 66812 147812 66876
rect 147876 66874 147882 66876
rect 333881 66874 333947 66877
rect 147876 66872 333947 66874
rect 147876 66816 333886 66872
rect 333942 66816 333947 66872
rect 147876 66814 333947 66816
rect 147876 66812 147882 66814
rect 333881 66811 333947 66814
rect 149973 65650 150039 65653
rect 149470 65648 150039 65650
rect 149470 65592 149978 65648
rect 150034 65592 150039 65648
rect 149470 65590 150039 65592
rect 149237 65378 149303 65381
rect 149470 65378 149530 65590
rect 149973 65587 150039 65590
rect 162710 65452 162716 65516
rect 162780 65514 162786 65516
rect 526621 65514 526687 65517
rect 162780 65512 526687 65514
rect 162780 65456 526626 65512
rect 526682 65456 526687 65512
rect 162780 65454 526687 65456
rect 162780 65452 162786 65454
rect 526621 65451 526687 65454
rect 149237 65376 149530 65378
rect 149237 65320 149242 65376
rect 149298 65320 149530 65376
rect 149237 65318 149530 65320
rect 149237 65315 149303 65318
rect 143390 64228 143396 64292
rect 143460 64290 143466 64292
rect 279509 64290 279575 64293
rect 143460 64288 279575 64290
rect 143460 64232 279514 64288
rect 279570 64232 279575 64288
rect 143460 64230 279575 64232
rect 143460 64228 143466 64230
rect 279509 64227 279575 64230
rect 52545 64154 52611 64157
rect 125726 64154 125732 64156
rect 52545 64152 125732 64154
rect 52545 64096 52550 64152
rect 52606 64096 125732 64152
rect 52545 64094 125732 64096
rect 52545 64091 52611 64094
rect 125726 64092 125732 64094
rect 125796 64092 125802 64156
rect 134742 64092 134748 64156
rect 134812 64154 134818 64156
rect 175457 64154 175523 64157
rect 134812 64152 175523 64154
rect 134812 64096 175462 64152
rect 175518 64096 175523 64152
rect 134812 64094 175523 64096
rect 134812 64092 134818 64094
rect 175457 64091 175523 64094
rect 178861 64154 178927 64157
rect 576117 64154 576183 64157
rect 178861 64152 576183 64154
rect 178861 64096 178866 64152
rect 178922 64096 576122 64152
rect 576178 64096 576183 64152
rect 178861 64094 576183 64096
rect 178861 64091 178927 64094
rect 576117 64091 576183 64094
rect 134926 62732 134932 62796
rect 134996 62794 135002 62796
rect 171961 62794 172027 62797
rect 134996 62792 172027 62794
rect 134996 62736 171966 62792
rect 172022 62736 172027 62792
rect 134996 62734 172027 62736
rect 134996 62732 135002 62734
rect 171961 62731 172027 62734
rect 87965 61434 88031 61437
rect 128670 61434 128676 61436
rect 87965 61432 128676 61434
rect 87965 61376 87970 61432
rect 88026 61376 128676 61432
rect 87965 61374 128676 61376
rect 87965 61371 88031 61374
rect 128670 61372 128676 61374
rect 128740 61372 128746 61436
rect 136030 61372 136036 61436
rect 136100 61434 136106 61436
rect 189717 61434 189783 61437
rect 136100 61432 189783 61434
rect 136100 61376 189722 61432
rect 189778 61376 189783 61432
rect 136100 61374 189783 61376
rect 136100 61372 136106 61374
rect 189717 61371 189783 61374
rect 155166 59876 155172 59940
rect 155236 59938 155242 59940
rect 439129 59938 439195 59941
rect 155236 59936 439195 59938
rect 155236 59880 439134 59936
rect 439190 59880 439195 59936
rect 155236 59878 439195 59880
rect 155236 59876 155242 59878
rect 439129 59875 439195 59878
rect 114369 59666 114435 59669
rect 583520 59666 584960 59756
rect 114369 59664 584960 59666
rect 114369 59608 114374 59664
rect 114430 59608 584960 59664
rect 114369 59606 584960 59608
rect 114369 59603 114435 59606
rect 583520 59516 584960 59606
rect 70301 58714 70367 58717
rect 127382 58714 127388 58716
rect 70301 58712 127388 58714
rect -960 58578 480 58668
rect 70301 58656 70306 58712
rect 70362 58656 127388 58712
rect 70301 58654 127388 58656
rect 70301 58651 70367 58654
rect 127382 58652 127388 58654
rect 127452 58652 127458 58716
rect 145046 58652 145052 58716
rect 145116 58714 145122 58716
rect 317321 58714 317387 58717
rect 145116 58712 317387 58714
rect 145116 58656 317326 58712
rect 317382 58656 317387 58712
rect 145116 58654 317387 58656
rect 145116 58652 145122 58654
rect 317321 58651 317387 58654
rect 3693 58578 3759 58581
rect -960 58576 3759 58578
rect -960 58520 3698 58576
rect 3754 58520 3759 58576
rect -960 58518 3759 58520
rect -960 58428 480 58518
rect 3693 58515 3759 58518
rect 114461 58578 114527 58581
rect 472617 58578 472683 58581
rect 114461 58576 472683 58578
rect 114461 58520 114466 58576
rect 114522 58520 472622 58576
rect 472678 58520 472683 58576
rect 114461 58518 472683 58520
rect 114461 58515 114527 58518
rect 472617 58515 472683 58518
rect 136214 57428 136220 57492
rect 136284 57490 136290 57492
rect 193213 57490 193279 57493
rect 136284 57488 193279 57490
rect 136284 57432 193218 57488
rect 193274 57432 193279 57488
rect 136284 57430 193279 57432
rect 136284 57428 136290 57430
rect 193213 57427 193279 57430
rect 157742 57292 157748 57356
rect 157812 57354 157818 57356
rect 474549 57354 474615 57357
rect 157812 57352 474615 57354
rect 157812 57296 474554 57352
rect 474610 57296 474615 57352
rect 157812 57294 474615 57296
rect 157812 57292 157818 57294
rect 474549 57291 474615 57294
rect 162342 57156 162348 57220
rect 162412 57218 162418 57220
rect 530117 57218 530183 57221
rect 162412 57216 530183 57218
rect 162412 57160 530122 57216
rect 530178 57160 530183 57216
rect 162412 57158 530183 57160
rect 162412 57156 162418 57158
rect 530117 57155 530183 57158
rect 137318 55932 137324 55996
rect 137388 55994 137394 55996
rect 210969 55994 211035 55997
rect 137388 55992 211035 55994
rect 137388 55936 210974 55992
rect 211030 55936 211035 55992
rect 137388 55934 211035 55936
rect 137388 55932 137394 55934
rect 210969 55931 211035 55934
rect 91553 55858 91619 55861
rect 128486 55858 128492 55860
rect 91553 55856 128492 55858
rect 91553 55800 91558 55856
rect 91614 55800 128492 55856
rect 91553 55798 128492 55800
rect 91553 55795 91619 55798
rect 128486 55796 128492 55798
rect 128556 55796 128562 55860
rect 161054 55796 161060 55860
rect 161124 55858 161130 55860
rect 512453 55858 512519 55861
rect 161124 55856 512519 55858
rect 161124 55800 512458 55856
rect 512514 55800 512519 55856
rect 161124 55798 512519 55800
rect 161124 55796 161130 55798
rect 512453 55795 512519 55798
rect 140078 54572 140084 54636
rect 140148 54634 140154 54636
rect 242893 54634 242959 54637
rect 140148 54632 242959 54634
rect 140148 54576 242898 54632
rect 242954 54576 242959 54632
rect 140148 54574 242959 54576
rect 140148 54572 140154 54574
rect 242893 54571 242959 54574
rect 159214 54436 159220 54500
rect 159284 54498 159290 54500
rect 494697 54498 494763 54501
rect 159284 54496 494763 54498
rect 159284 54440 494702 54496
rect 494758 54440 494763 54496
rect 159284 54438 494763 54440
rect 159284 54436 159290 54438
rect 494697 54435 494763 54438
rect 38377 53138 38443 53141
rect 124622 53138 124628 53140
rect 38377 53136 124628 53138
rect 38377 53080 38382 53136
rect 38438 53080 124628 53136
rect 38377 53078 124628 53080
rect 38377 53075 38443 53078
rect 124622 53076 124628 53078
rect 124692 53076 124698 53140
rect 135110 51988 135116 52052
rect 135180 52050 135186 52052
rect 174261 52050 174327 52053
rect 135180 52048 174327 52050
rect 135180 51992 174266 52048
rect 174322 51992 174327 52048
rect 135180 51990 174327 51992
rect 135180 51988 135186 51990
rect 174261 51987 174327 51990
rect 140262 51852 140268 51916
rect 140332 51914 140338 51916
rect 246389 51914 246455 51917
rect 140332 51912 246455 51914
rect 140332 51856 246394 51912
rect 246450 51856 246455 51912
rect 140332 51854 246455 51856
rect 140332 51852 140338 51854
rect 246389 51851 246455 51854
rect 18597 51778 18663 51781
rect 123334 51778 123340 51780
rect 18597 51776 123340 51778
rect 18597 51720 18602 51776
rect 18658 51720 123340 51776
rect 18597 51718 123340 51720
rect 18597 51715 18663 51718
rect 123334 51716 123340 51718
rect 123404 51716 123410 51780
rect 155350 51716 155356 51780
rect 155420 51778 155426 51780
rect 437933 51778 437999 51781
rect 155420 51776 437999 51778
rect 155420 51720 437938 51776
rect 437994 51720 437999 51776
rect 155420 51718 437999 51720
rect 155420 51716 155426 51718
rect 437933 51715 437999 51718
rect 73797 50418 73863 50421
rect 127198 50418 127204 50420
rect 73797 50416 127204 50418
rect 73797 50360 73802 50416
rect 73858 50360 127204 50416
rect 73797 50358 127204 50360
rect 73797 50355 73863 50358
rect 127198 50356 127204 50358
rect 127268 50356 127274 50420
rect 143022 50356 143028 50420
rect 143092 50418 143098 50420
rect 278313 50418 278379 50421
rect 143092 50416 278379 50418
rect 143092 50360 278318 50416
rect 278374 50360 278379 50416
rect 143092 50358 278379 50360
rect 143092 50356 143098 50358
rect 278313 50355 278379 50358
rect 40769 50282 40835 50285
rect 124438 50282 124444 50284
rect 40769 50280 124444 50282
rect 40769 50224 40774 50280
rect 40830 50224 124444 50280
rect 40769 50222 124444 50224
rect 40769 50219 40835 50222
rect 124438 50220 124444 50222
rect 124508 50220 124514 50284
rect 161238 50220 161244 50284
rect 161308 50282 161314 50284
rect 511257 50282 511323 50285
rect 161308 50280 511323 50282
rect 161308 50224 511262 50280
rect 511318 50224 511323 50280
rect 161308 50222 511323 50224
rect 161308 50220 161314 50222
rect 511257 50219 511323 50222
rect 74993 49058 75059 49061
rect 127014 49058 127020 49060
rect 74993 49056 127020 49058
rect 74993 49000 74998 49056
rect 75054 49000 127020 49056
rect 74993 48998 127020 49000
rect 74993 48995 75059 48998
rect 127014 48996 127020 48998
rect 127084 48996 127090 49060
rect 143206 48996 143212 49060
rect 143276 49058 143282 49060
rect 281901 49058 281967 49061
rect 143276 49056 281967 49058
rect 143276 49000 281906 49056
rect 281962 49000 281967 49056
rect 143276 48998 281967 49000
rect 143276 48996 143282 48998
rect 281901 48995 281967 48998
rect 37917 48922 37983 48925
rect 124806 48922 124812 48924
rect 37917 48920 124812 48922
rect 37917 48864 37922 48920
rect 37978 48864 124812 48920
rect 37917 48862 124812 48864
rect 37917 48859 37983 48862
rect 124806 48860 124812 48862
rect 124876 48860 124882 48924
rect 165102 48860 165108 48924
rect 165172 48922 165178 48924
rect 565629 48922 565695 48925
rect 165172 48920 565695 48922
rect 165172 48864 565634 48920
rect 565690 48864 565695 48920
rect 165172 48862 565695 48864
rect 165172 48860 165178 48862
rect 565629 48859 565695 48862
rect 133086 48180 133092 48244
rect 133156 48242 133162 48244
rect 136265 48242 136331 48245
rect 133156 48240 136331 48242
rect 133156 48184 136270 48240
rect 136326 48184 136331 48240
rect 133156 48182 136331 48184
rect 133156 48180 133162 48182
rect 136265 48179 136331 48182
rect 147070 47636 147076 47700
rect 147140 47698 147146 47700
rect 331581 47698 331647 47701
rect 147140 47696 331647 47698
rect 147140 47640 331586 47696
rect 331642 47640 331647 47696
rect 147140 47638 331647 47640
rect 147140 47636 147146 47638
rect 331581 47635 331647 47638
rect 166390 47500 166396 47564
rect 166460 47562 166466 47564
rect 576301 47562 576367 47565
rect 166460 47560 576367 47562
rect 166460 47504 576306 47560
rect 576362 47504 576367 47560
rect 166460 47502 576367 47504
rect 166460 47500 166466 47502
rect 576301 47499 576367 47502
rect 147254 46548 147260 46612
rect 147324 46610 147330 46612
rect 335077 46610 335143 46613
rect 147324 46608 335143 46610
rect 147324 46552 335082 46608
rect 335138 46552 335143 46608
rect 147324 46550 335143 46552
rect 147324 46548 147330 46550
rect 335077 46547 335143 46550
rect 151118 46412 151124 46476
rect 151188 46474 151194 46476
rect 384757 46474 384823 46477
rect 151188 46472 384823 46474
rect 151188 46416 384762 46472
rect 384818 46416 384823 46472
rect 151188 46414 384823 46416
rect 151188 46412 151194 46414
rect 384757 46411 384823 46414
rect 178769 46338 178835 46341
rect 583520 46338 584960 46428
rect 178769 46336 584960 46338
rect 178769 46280 178774 46336
rect 178830 46280 584960 46336
rect 178769 46278 584960 46280
rect 178769 46275 178835 46278
rect 53741 46202 53807 46205
rect 125542 46202 125548 46204
rect 53741 46200 125548 46202
rect 53741 46144 53746 46200
rect 53802 46144 125548 46200
rect 53741 46142 125548 46144
rect 53741 46139 53807 46142
rect 125542 46140 125548 46142
rect 125612 46140 125618 46204
rect 167494 46140 167500 46204
rect 167564 46202 167570 46204
rect 580993 46202 581059 46205
rect 167564 46200 581059 46202
rect 167564 46144 580998 46200
rect 581054 46144 581059 46200
rect 583520 46188 584960 46278
rect 167564 46142 581059 46144
rect 167564 46140 167570 46142
rect 580993 46139 581059 46142
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 147990 44780 147996 44844
rect 148060 44842 148066 44844
rect 349245 44842 349311 44845
rect 148060 44840 349311 44842
rect 148060 44784 349250 44840
rect 349306 44784 349311 44840
rect 148060 44782 349311 44784
rect 148060 44780 148066 44782
rect 349245 44779 349311 44782
rect 148174 43420 148180 43484
rect 148244 43482 148250 43484
rect 352833 43482 352899 43485
rect 148244 43480 352899 43482
rect 148244 43424 352838 43480
rect 352894 43424 352899 43480
rect 148244 43422 352899 43424
rect 148244 43420 148250 43422
rect 352833 43419 352899 43422
rect 133270 42060 133276 42124
rect 133340 42122 133346 42124
rect 156597 42122 156663 42125
rect 133340 42120 156663 42122
rect 133340 42064 156602 42120
rect 156658 42064 156663 42120
rect 133340 42062 156663 42064
rect 133340 42060 133346 42062
rect 156597 42059 156663 42062
rect 163446 42060 163452 42124
rect 163516 42122 163522 42124
rect 547873 42122 547939 42125
rect 163516 42120 547939 42122
rect 163516 42064 547878 42120
rect 547934 42064 547939 42120
rect 163516 42062 547939 42064
rect 163516 42060 163522 42062
rect 547873 42059 547939 42062
rect 150198 40700 150204 40764
rect 150268 40762 150274 40764
rect 370589 40762 370655 40765
rect 150268 40760 370655 40762
rect 150268 40704 370594 40760
rect 370650 40704 370655 40760
rect 150268 40702 370655 40704
rect 150268 40700 150274 40702
rect 370589 40699 370655 40702
rect 153878 40564 153884 40628
rect 153948 40626 153954 40628
rect 420177 40626 420243 40629
rect 153948 40624 420243 40626
rect 153948 40568 420182 40624
rect 420238 40568 420243 40624
rect 153948 40566 420243 40568
rect 153948 40564 153954 40566
rect 420177 40563 420243 40566
rect 136398 39340 136404 39404
rect 136468 39402 136474 39404
rect 190821 39402 190887 39405
rect 136468 39400 190887 39402
rect 136468 39344 190826 39400
rect 190882 39344 190887 39400
rect 136468 39342 190887 39344
rect 136468 39340 136474 39342
rect 190821 39339 190887 39342
rect 151302 39204 151308 39268
rect 151372 39266 151378 39268
rect 388253 39266 388319 39269
rect 151372 39264 388319 39266
rect 151372 39208 388258 39264
rect 388314 39208 388319 39264
rect 151372 39206 388319 39208
rect 151372 39204 151378 39206
rect 388253 39203 388319 39206
rect 133454 37980 133460 38044
rect 133524 38042 133530 38044
rect 155217 38042 155283 38045
rect 133524 38040 155283 38042
rect 133524 37984 155222 38040
rect 155278 37984 155283 38040
rect 133524 37982 155283 37984
rect 133524 37980 133530 37982
rect 155217 37979 155283 37982
rect 152222 37844 152228 37908
rect 152292 37906 152298 37908
rect 406009 37906 406075 37909
rect 152292 37904 406075 37906
rect 152292 37848 406014 37904
rect 406070 37848 406075 37904
rect 152292 37846 406075 37848
rect 152292 37844 152298 37846
rect 406009 37843 406075 37846
rect 140446 36620 140452 36684
rect 140516 36682 140522 36684
rect 244089 36682 244155 36685
rect 140516 36680 244155 36682
rect 140516 36624 244094 36680
rect 244150 36624 244155 36680
rect 140516 36622 244155 36624
rect 140516 36620 140522 36622
rect 244089 36619 244155 36622
rect 154062 36484 154068 36548
rect 154132 36546 154138 36548
rect 423765 36546 423831 36549
rect 154132 36544 423831 36546
rect 154132 36488 423770 36544
rect 423826 36488 423831 36544
rect 154132 36486 423831 36488
rect 154132 36484 154138 36486
rect 423765 36483 423831 36486
rect 155534 35260 155540 35324
rect 155604 35322 155610 35324
rect 441521 35322 441587 35325
rect 155604 35320 441587 35322
rect 155604 35264 441526 35320
rect 441582 35264 441587 35320
rect 155604 35262 441587 35264
rect 155604 35260 155610 35262
rect 441521 35259 441587 35262
rect 156086 35124 156092 35188
rect 156156 35186 156162 35188
rect 456885 35186 456951 35189
rect 156156 35184 456951 35186
rect 156156 35128 456890 35184
rect 456946 35128 456951 35184
rect 156156 35126 456951 35128
rect 156156 35124 156162 35126
rect 456885 35123 456951 35126
rect 3417 33962 3483 33965
rect 177021 33962 177087 33965
rect 3417 33960 177087 33962
rect 3417 33904 3422 33960
rect 3478 33904 177026 33960
rect 177082 33904 177087 33960
rect 3417 33902 177087 33904
rect 3417 33899 3483 33902
rect 177021 33899 177087 33902
rect 151486 33764 151492 33828
rect 151556 33826 151562 33828
rect 387149 33826 387215 33829
rect 151556 33824 387215 33826
rect 151556 33768 387154 33824
rect 387210 33768 387215 33824
rect 151556 33766 387215 33768
rect 151556 33764 151562 33766
rect 387149 33763 387215 33766
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 155718 30908 155724 30972
rect 155788 30970 155794 30972
rect 440325 30970 440391 30973
rect 155788 30968 440391 30970
rect 155788 30912 440330 30968
rect 440386 30912 440391 30968
rect 155788 30910 440391 30912
rect 155788 30908 155794 30910
rect 440325 30907 440391 30910
rect 165286 29548 165292 29612
rect 165356 29610 165362 29612
rect 563237 29610 563303 29613
rect 165356 29608 563303 29610
rect 165356 29552 563242 29608
rect 563298 29552 563303 29608
rect 165356 29550 563303 29552
rect 165356 29548 165362 29550
rect 563237 29547 563303 29550
rect 137502 26964 137508 27028
rect 137572 27026 137578 27028
rect 209773 27026 209839 27029
rect 137572 27024 209839 27026
rect 137572 26968 209778 27024
rect 209834 26968 209839 27024
rect 137572 26966 209839 26968
rect 137572 26964 137578 26966
rect 209773 26963 209839 26966
rect 159398 26828 159404 26892
rect 159468 26890 159474 26892
rect 492305 26890 492371 26893
rect 159468 26888 492371 26890
rect 159468 26832 492310 26888
rect 492366 26832 492371 26888
rect 159468 26830 492371 26832
rect 159468 26828 159474 26830
rect 492305 26827 492371 26830
rect 139158 25604 139164 25668
rect 139228 25666 139234 25668
rect 226333 25666 226399 25669
rect 139228 25664 226399 25666
rect 139228 25608 226338 25664
rect 226394 25608 226399 25664
rect 139228 25606 226399 25608
rect 139228 25604 139234 25606
rect 226333 25603 226399 25606
rect 152406 25468 152412 25532
rect 152476 25530 152482 25532
rect 404813 25530 404879 25533
rect 152476 25528 404879 25530
rect 152476 25472 404818 25528
rect 404874 25472 404879 25528
rect 152476 25470 404879 25472
rect 152476 25468 152482 25470
rect 404813 25467 404879 25470
rect 146886 22748 146892 22812
rect 146956 22810 146962 22812
rect 332685 22810 332751 22813
rect 146956 22808 332751 22810
rect 146956 22752 332690 22808
rect 332746 22752 332751 22808
rect 146956 22750 332751 22752
rect 146956 22748 146962 22750
rect 332685 22747 332751 22750
rect 154246 22612 154252 22676
rect 154316 22674 154322 22676
rect 421373 22674 421439 22677
rect 154316 22672 421439 22674
rect 154316 22616 421378 22672
rect 421434 22616 421439 22672
rect 154316 22614 421439 22616
rect 154316 22612 154322 22614
rect 421373 22611 421439 22614
rect 148358 21252 148364 21316
rect 148428 21314 148434 21316
rect 351637 21314 351703 21317
rect 148428 21312 351703 21314
rect 148428 21256 351642 21312
rect 351698 21256 351703 21312
rect 148428 21254 351703 21256
rect 148428 21252 148434 21254
rect 351637 21251 351703 21254
rect 142838 19892 142844 19956
rect 142908 19954 142914 19956
rect 280705 19954 280771 19957
rect 142908 19952 280771 19954
rect 142908 19896 280710 19952
rect 280766 19896 280771 19952
rect 142908 19894 280771 19896
rect 142908 19892 142914 19894
rect 280705 19891 280771 19894
rect 472617 19818 472683 19821
rect 583520 19818 584960 19908
rect 472617 19816 584960 19818
rect 472617 19760 472622 19816
rect 472678 19760 584960 19816
rect 472617 19758 584960 19760
rect 472617 19755 472683 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3601 19410 3667 19413
rect -960 19408 3667 19410
rect -960 19352 3606 19408
rect 3662 19352 3667 19408
rect -960 19350 3667 19352
rect -960 19260 480 19350
rect 3601 19347 3667 19350
rect 165470 18668 165476 18732
rect 165540 18730 165546 18732
rect 564433 18730 564499 18733
rect 165540 18728 564499 18730
rect 165540 18672 564438 18728
rect 564494 18672 564499 18728
rect 165540 18670 564499 18672
rect 165540 18668 165546 18670
rect 564433 18667 564499 18670
rect 166574 18532 166580 18596
rect 166644 18594 166650 18596
rect 578601 18594 578667 18597
rect 166644 18592 578667 18594
rect 166644 18536 578606 18592
rect 578662 18536 578667 18592
rect 166644 18534 578667 18536
rect 166644 18532 166650 18534
rect 578601 18531 578667 18534
rect 131982 17172 131988 17236
rect 132052 17234 132058 17236
rect 140037 17234 140103 17237
rect 132052 17232 140103 17234
rect 132052 17176 140042 17232
rect 140098 17176 140103 17232
rect 132052 17174 140103 17176
rect 132052 17172 132058 17174
rect 140037 17171 140103 17174
rect 133638 15812 133644 15876
rect 133708 15874 133714 15876
rect 151169 15874 151235 15877
rect 133708 15872 151235 15874
rect 133708 15816 151174 15872
rect 151230 15816 151235 15872
rect 133708 15814 151235 15816
rect 133708 15812 133714 15814
rect 151169 15811 151235 15814
rect 159582 15812 159588 15876
rect 159652 15874 159658 15876
rect 489913 15874 489979 15877
rect 159652 15872 489979 15874
rect 159652 15816 489918 15872
rect 489974 15816 489979 15872
rect 159652 15814 489979 15816
rect 159652 15812 159658 15814
rect 489913 15811 489979 15814
rect 162526 14452 162532 14516
rect 162596 14514 162602 14516
rect 529013 14514 529079 14517
rect 162596 14512 529079 14514
rect 162596 14456 529018 14512
rect 529074 14456 529079 14512
rect 162596 14454 529079 14456
rect 162596 14452 162602 14454
rect 529013 14451 529079 14454
rect 166758 12956 166764 13020
rect 166828 13018 166834 13020
rect 577405 13018 577471 13021
rect 166828 13016 577471 13018
rect 166828 12960 577410 13016
rect 577466 12960 577471 13016
rect 166828 12958 577471 12960
rect 166828 12956 166834 12958
rect 577405 12955 577471 12958
rect 140630 11868 140636 11932
rect 140700 11930 140706 11932
rect 245193 11930 245259 11933
rect 140700 11928 245259 11930
rect 140700 11872 245198 11928
rect 245254 11872 245259 11928
rect 140700 11870 245259 11872
rect 140700 11868 140706 11870
rect 245193 11867 245259 11870
rect 151670 11732 151676 11796
rect 151740 11794 151746 11796
rect 385953 11794 386019 11797
rect 151740 11792 386019 11794
rect 151740 11736 385958 11792
rect 386014 11736 386019 11792
rect 151740 11734 386019 11736
rect 151740 11732 151746 11734
rect 385953 11731 386019 11734
rect 162158 11596 162164 11660
rect 162228 11658 162234 11660
rect 527817 11658 527883 11661
rect 162228 11656 527883 11658
rect 162228 11600 527822 11656
rect 527878 11600 527883 11656
rect 162228 11598 527883 11600
rect 162228 11596 162234 11598
rect 527817 11595 527883 11598
rect 148542 10236 148548 10300
rect 148612 10298 148618 10300
rect 350441 10298 350507 10301
rect 148612 10296 350507 10298
rect 148612 10240 350446 10296
rect 350502 10240 350507 10296
rect 148612 10238 350507 10240
rect 148612 10236 148618 10238
rect 350441 10235 350507 10238
rect 144310 9012 144316 9076
rect 144380 9074 144386 9076
rect 297265 9074 297331 9077
rect 144380 9072 297331 9074
rect 144380 9016 297270 9072
rect 297326 9016 297331 9072
rect 144380 9014 297331 9016
rect 144380 9012 144386 9014
rect 297265 9011 297331 9014
rect 146150 8876 146156 8940
rect 146220 8938 146226 8940
rect 316217 8938 316283 8941
rect 146220 8936 316283 8938
rect 146220 8880 316222 8936
rect 316278 8880 316283 8936
rect 146220 8878 316283 8880
rect 146220 8876 146226 8878
rect 316217 8875 316283 8878
rect 154430 7516 154436 7580
rect 154500 7578 154506 7580
rect 418981 7578 419047 7581
rect 154500 7576 419047 7578
rect 154500 7520 418986 7576
rect 419042 7520 419047 7576
rect 154500 7518 419047 7520
rect 154500 7516 154506 7518
rect 418981 7515 419047 7518
rect 576117 6626 576183 6629
rect 583520 6626 584960 6716
rect 576117 6624 584960 6626
rect -960 6490 480 6580
rect 576117 6568 576122 6624
rect 576178 6568 584960 6624
rect 576117 6566 584960 6568
rect 576117 6563 576183 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 132166 6428 132172 6492
rect 132236 6490 132242 6492
rect 255865 6490 255931 6493
rect 132236 6488 255931 6490
rect 132236 6432 255870 6488
rect 255926 6432 255931 6488
rect 583520 6476 584960 6566
rect 132236 6430 255931 6432
rect 132236 6428 132242 6430
rect 255865 6427 255931 6430
rect 158294 6292 158300 6356
rect 158364 6354 158370 6356
rect 473445 6354 473511 6357
rect 158364 6352 473511 6354
rect 158364 6296 473450 6352
rect 473506 6296 473511 6352
rect 158364 6294 473511 6296
rect 158364 6292 158370 6294
rect 473445 6291 473511 6294
rect 89161 6218 89227 6221
rect 128854 6218 128860 6220
rect 89161 6216 128860 6218
rect 89161 6160 89166 6216
rect 89222 6160 128860 6216
rect 89161 6158 128860 6160
rect 89161 6155 89227 6158
rect 128854 6156 128860 6158
rect 128924 6156 128930 6220
rect 157926 6156 157932 6220
rect 157996 6218 158002 6220
rect 476941 6218 477007 6221
rect 157996 6216 477007 6218
rect 157996 6160 476946 6216
rect 477002 6160 477007 6216
rect 157996 6158 477007 6160
rect 157996 6156 158002 6158
rect 476941 6155 477007 6158
rect 159766 4796 159772 4860
rect 159836 4858 159842 4860
rect 493501 4858 493567 4861
rect 159836 4856 493567 4858
rect 159836 4800 493506 4856
rect 493562 4800 493567 4856
rect 159836 4798 493567 4800
rect 159836 4796 159842 4798
rect 493501 4795 493567 4798
rect 130878 3844 130884 3908
rect 130948 3906 130954 3908
rect 161289 3906 161355 3909
rect 130948 3904 161355 3906
rect 130948 3848 161294 3904
rect 161350 3848 161355 3904
rect 130948 3846 161355 3848
rect 130948 3844 130954 3846
rect 161289 3843 161355 3846
rect 141182 3708 141188 3772
rect 141252 3770 141258 3772
rect 264145 3770 264211 3773
rect 141252 3768 264211 3770
rect 141252 3712 264150 3768
rect 264206 3712 264211 3768
rect 141252 3710 264211 3712
rect 141252 3708 141258 3710
rect 264145 3707 264211 3710
rect 144126 3572 144132 3636
rect 144196 3634 144202 3636
rect 296069 3634 296135 3637
rect 144196 3632 296135 3634
rect 144196 3576 296074 3632
rect 296130 3576 296135 3632
rect 144196 3574 296135 3576
rect 144196 3572 144202 3574
rect 296069 3571 296135 3574
rect 144494 3436 144500 3500
rect 144564 3498 144570 3500
rect 299657 3498 299723 3501
rect 144564 3496 299723 3498
rect 144564 3440 299662 3496
rect 299718 3440 299723 3496
rect 144564 3438 299723 3440
rect 144564 3436 144570 3438
rect 299657 3435 299723 3438
rect 132350 3300 132356 3364
rect 132420 3362 132426 3364
rect 138841 3362 138907 3365
rect 132420 3360 138907 3362
rect 132420 3304 138846 3360
rect 138902 3304 138907 3360
rect 132420 3302 138907 3304
rect 132420 3300 132426 3302
rect 138841 3299 138907 3302
rect 157190 3300 157196 3364
rect 157260 3362 157266 3364
rect 459185 3362 459251 3365
rect 157260 3360 459251 3362
rect 157260 3304 459190 3360
rect 459246 3304 459251 3360
rect 157260 3302 459251 3304
rect 157260 3300 157266 3302
rect 459185 3299 459251 3302
<< via3 >>
rect 136036 181052 136100 181116
rect 135852 180916 135916 180980
rect 140636 178068 140700 178132
rect 139532 177380 139596 177444
rect 141924 176020 141988 176084
rect 141556 172484 141620 172548
rect 139532 165200 139596 165204
rect 139532 165144 139546 165200
rect 139546 165144 139596 165200
rect 139532 165140 139596 165144
rect 141556 162148 141620 162212
rect 135852 161468 135916 161532
rect 136404 161332 136468 161396
rect 135852 159972 135916 160036
rect 136036 159972 136100 160036
rect 140636 152356 140700 152420
rect 135852 137532 135916 137596
rect 136036 137396 136100 137460
rect 141924 137396 141988 137460
rect 169340 75380 169404 75444
rect 147444 75244 147508 75308
rect 160876 75108 160940 75172
rect 158852 74836 158916 74900
rect 161428 74836 161492 74900
rect 155908 74700 155972 74764
rect 157196 74564 157260 74628
rect 169340 74564 169404 74628
rect 151492 73884 151556 73948
rect 157196 73884 157260 73948
rect 140268 73612 140332 73676
rect 123708 73536 123772 73540
rect 123708 73480 123722 73536
rect 123722 73480 123772 73536
rect 123708 73476 123772 73480
rect 139164 73536 139228 73540
rect 139164 73480 139178 73536
rect 139178 73480 139228 73536
rect 139164 73476 139228 73480
rect 140452 73536 140516 73540
rect 140452 73480 140502 73536
rect 140502 73480 140516 73536
rect 140452 73476 140516 73480
rect 141188 73476 141252 73540
rect 139348 73340 139412 73404
rect 140084 73340 140148 73404
rect 140636 73400 140700 73404
rect 140636 73344 140650 73400
rect 140650 73344 140700 73400
rect 140636 73340 140700 73344
rect 158852 73400 158916 73404
rect 161612 73476 161676 73540
rect 166212 73476 166276 73540
rect 158852 73344 158902 73400
rect 158902 73344 158916 73400
rect 158852 73340 158916 73344
rect 161244 73264 161308 73268
rect 161244 73208 161294 73264
rect 161294 73208 161308 73264
rect 161244 73204 161308 73208
rect 147444 73068 147508 73132
rect 147996 73068 148060 73132
rect 124444 72796 124508 72860
rect 125548 72796 125612 72860
rect 121500 72660 121564 72724
rect 123156 72720 123220 72724
rect 123156 72664 123206 72720
rect 123206 72664 123220 72720
rect 123156 72660 123220 72664
rect 124260 72720 124324 72724
rect 124260 72664 124274 72720
rect 124274 72664 124324 72720
rect 124260 72660 124324 72664
rect 124628 72660 124692 72724
rect 125732 72660 125796 72724
rect 123708 72584 123772 72588
rect 123708 72528 123758 72584
rect 123758 72528 123772 72584
rect 123708 72524 123772 72528
rect 124812 72524 124876 72588
rect 127388 72796 127452 72860
rect 128676 72796 128740 72860
rect 130884 72932 130948 72996
rect 142844 72932 142908 72996
rect 131988 72796 132052 72860
rect 133276 72796 133340 72860
rect 135116 72856 135180 72860
rect 135116 72800 135130 72856
rect 135130 72800 135180 72856
rect 135116 72796 135180 72800
rect 136588 72796 136652 72860
rect 137324 72796 137388 72860
rect 143396 72796 143460 72860
rect 144500 72796 144564 72860
rect 145052 72796 145116 72860
rect 147628 72932 147692 72996
rect 148364 72796 148428 72860
rect 150388 72796 150452 72860
rect 152228 72796 152292 72860
rect 153884 72796 153948 72860
rect 155356 72796 155420 72860
rect 127204 72720 127268 72724
rect 127204 72664 127254 72720
rect 127254 72664 127268 72720
rect 127204 72660 127268 72664
rect 128492 72660 128556 72724
rect 132356 72720 132420 72724
rect 132356 72664 132370 72720
rect 132370 72664 132420 72720
rect 132356 72660 132420 72664
rect 133644 72720 133708 72724
rect 133644 72664 133658 72720
rect 133658 72664 133708 72720
rect 133644 72660 133708 72664
rect 134932 72720 134996 72724
rect 134932 72664 134946 72720
rect 134946 72664 134996 72720
rect 134932 72660 134996 72664
rect 136404 72720 136468 72724
rect 136404 72664 136418 72720
rect 136418 72664 136468 72720
rect 136404 72660 136468 72664
rect 137508 72660 137572 72724
rect 143028 72660 143092 72724
rect 144868 72660 144932 72724
rect 146156 72720 146220 72724
rect 146156 72664 146170 72720
rect 146170 72664 146220 72720
rect 146156 72660 146220 72664
rect 147076 72660 147140 72724
rect 127572 72524 127636 72588
rect 128860 72524 128924 72588
rect 133092 72524 133156 72588
rect 134748 72524 134812 72588
rect 136220 72524 136284 72588
rect 143212 72524 143276 72588
rect 144316 72524 144380 72588
rect 123340 72388 123404 72452
rect 127020 72388 127084 72452
rect 133460 72388 133524 72452
rect 134564 72388 134628 72452
rect 136036 72388 136100 72452
rect 132172 72252 132236 72316
rect 144132 72388 144196 72452
rect 148548 72660 148612 72724
rect 150204 72660 150268 72724
rect 151676 72660 151740 72724
rect 152412 72660 152476 72724
rect 154252 72720 154316 72724
rect 154252 72664 154302 72720
rect 154302 72664 154316 72720
rect 154252 72660 154316 72664
rect 155724 72720 155788 72724
rect 155724 72664 155774 72720
rect 155774 72664 155788 72720
rect 155724 72660 155788 72664
rect 157564 73128 157628 73132
rect 157564 73072 157578 73128
rect 157578 73072 157628 73128
rect 157564 73068 157628 73072
rect 162164 73068 162228 73132
rect 159036 72932 159100 72996
rect 158300 72720 158364 72724
rect 158300 72664 158350 72720
rect 158350 72664 158364 72720
rect 158300 72660 158364 72664
rect 158668 72660 158732 72724
rect 159220 72720 159284 72724
rect 159220 72664 159234 72720
rect 159234 72664 159284 72720
rect 159220 72660 159284 72664
rect 159588 72720 159652 72724
rect 159588 72664 159638 72720
rect 159638 72664 159652 72720
rect 159588 72660 159652 72664
rect 159772 72660 159836 72724
rect 162532 72660 162596 72724
rect 163452 72660 163516 72724
rect 165292 72720 165356 72724
rect 165292 72664 165342 72720
rect 165342 72664 165356 72720
rect 165292 72660 165356 72664
rect 148180 72524 148244 72588
rect 151124 72524 151188 72588
rect 154068 72524 154132 72588
rect 155172 72524 155236 72588
rect 157196 72584 157260 72588
rect 157196 72528 157246 72584
rect 157246 72528 157260 72584
rect 157196 72524 157260 72528
rect 157932 72524 157996 72588
rect 159404 72524 159468 72588
rect 161060 72524 161124 72588
rect 162716 72524 162780 72588
rect 165476 72584 165540 72588
rect 165476 72528 165490 72584
rect 165490 72528 165540 72584
rect 165476 72524 165540 72528
rect 166580 72584 166644 72588
rect 166580 72528 166594 72584
rect 166594 72528 166644 72584
rect 166580 72524 166644 72528
rect 151308 72388 151372 72452
rect 154436 72388 154500 72452
rect 155540 72388 155604 72452
rect 146892 72116 146956 72180
rect 157748 72388 157812 72452
rect 159036 72388 159100 72452
rect 161428 72252 161492 72316
rect 162348 72388 162412 72452
rect 163084 72388 163148 72452
rect 165108 72388 165172 72452
rect 166764 72388 166828 72452
rect 157564 72116 157628 72180
rect 166396 72176 166460 72180
rect 166396 72120 166410 72176
rect 166410 72120 166460 72176
rect 166396 72116 166460 72120
rect 167500 72116 167564 72180
rect 160876 71980 160940 72044
rect 147628 71844 147692 71908
rect 155908 71844 155972 71908
rect 156092 71844 156156 71908
rect 166212 71844 166276 71908
rect 147444 71496 147508 71500
rect 147444 71440 147494 71496
rect 147494 71440 147508 71496
rect 147444 71436 147508 71440
rect 147260 71300 147324 71364
rect 161612 71300 161676 71364
rect 121500 69532 121564 69596
rect 150388 69532 150452 69596
rect 134564 68580 134628 68644
rect 136588 68444 136652 68508
rect 139348 68308 139412 68372
rect 127572 68172 127636 68236
rect 163084 68172 163148 68236
rect 158668 67084 158732 67148
rect 124260 66948 124324 67012
rect 144868 66948 144932 67012
rect 123156 66812 123220 66876
rect 147812 66812 147876 66876
rect 162716 65452 162780 65516
rect 143396 64228 143460 64292
rect 125732 64092 125796 64156
rect 134748 64092 134812 64156
rect 134932 62732 134996 62796
rect 128676 61372 128740 61436
rect 136036 61372 136100 61436
rect 155172 59876 155236 59940
rect 127388 58652 127452 58716
rect 145052 58652 145116 58716
rect 136220 57428 136284 57492
rect 157748 57292 157812 57356
rect 162348 57156 162412 57220
rect 137324 55932 137388 55996
rect 128492 55796 128556 55860
rect 161060 55796 161124 55860
rect 140084 54572 140148 54636
rect 159220 54436 159284 54500
rect 124628 53076 124692 53140
rect 135116 51988 135180 52052
rect 140268 51852 140332 51916
rect 123340 51716 123404 51780
rect 155356 51716 155420 51780
rect 127204 50356 127268 50420
rect 143028 50356 143092 50420
rect 124444 50220 124508 50284
rect 161244 50220 161308 50284
rect 127020 48996 127084 49060
rect 143212 48996 143276 49060
rect 124812 48860 124876 48924
rect 165108 48860 165172 48924
rect 133092 48180 133156 48244
rect 147076 47636 147140 47700
rect 166396 47500 166460 47564
rect 147260 46548 147324 46612
rect 151124 46412 151188 46476
rect 125548 46140 125612 46204
rect 167500 46140 167564 46204
rect 147996 44780 148060 44844
rect 148180 43420 148244 43484
rect 133276 42060 133340 42124
rect 163452 42060 163516 42124
rect 150204 40700 150268 40764
rect 153884 40564 153948 40628
rect 136404 39340 136468 39404
rect 151308 39204 151372 39268
rect 133460 37980 133524 38044
rect 152228 37844 152292 37908
rect 140452 36620 140516 36684
rect 154068 36484 154132 36548
rect 155540 35260 155604 35324
rect 156092 35124 156156 35188
rect 151492 33764 151556 33828
rect 155724 30908 155788 30972
rect 165292 29548 165356 29612
rect 137508 26964 137572 27028
rect 159404 26828 159468 26892
rect 139164 25604 139228 25668
rect 152412 25468 152476 25532
rect 146892 22748 146956 22812
rect 154252 22612 154316 22676
rect 148364 21252 148428 21316
rect 142844 19892 142908 19956
rect 165476 18668 165540 18732
rect 166580 18532 166644 18596
rect 131988 17172 132052 17236
rect 133644 15812 133708 15876
rect 159588 15812 159652 15876
rect 162532 14452 162596 14516
rect 166764 12956 166828 13020
rect 140636 11868 140700 11932
rect 151676 11732 151740 11796
rect 162164 11596 162228 11660
rect 148548 10236 148612 10300
rect 144316 9012 144380 9076
rect 146156 8876 146220 8940
rect 154436 7516 154500 7580
rect 132172 6428 132236 6492
rect 158300 6292 158364 6356
rect 128860 6156 128924 6220
rect 157932 6156 157996 6220
rect 159772 4796 159836 4860
rect 130884 3844 130948 3908
rect 141188 3708 141252 3772
rect 144132 3572 144196 3636
rect 144500 3436 144564 3500
rect 132356 3300 132420 3364
rect 157196 3300 157260 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 675494 -8106 711002
rect -8726 675258 -8694 675494
rect -8458 675258 -8374 675494
rect -8138 675258 -8106 675494
rect -8726 675174 -8106 675258
rect -8726 674938 -8694 675174
rect -8458 674938 -8374 675174
rect -8138 674938 -8106 675174
rect -8726 641494 -8106 674938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 607494 -8106 640938
rect -8726 607258 -8694 607494
rect -8458 607258 -8374 607494
rect -8138 607258 -8106 607494
rect -8726 607174 -8106 607258
rect -8726 606938 -8694 607174
rect -8458 606938 -8374 607174
rect -8138 606938 -8106 607174
rect -8726 573494 -8106 606938
rect -8726 573258 -8694 573494
rect -8458 573258 -8374 573494
rect -8138 573258 -8106 573494
rect -8726 573174 -8106 573258
rect -8726 572938 -8694 573174
rect -8458 572938 -8374 573174
rect -8138 572938 -8106 573174
rect -8726 539494 -8106 572938
rect -8726 539258 -8694 539494
rect -8458 539258 -8374 539494
rect -8138 539258 -8106 539494
rect -8726 539174 -8106 539258
rect -8726 538938 -8694 539174
rect -8458 538938 -8374 539174
rect -8138 538938 -8106 539174
rect -8726 505494 -8106 538938
rect -8726 505258 -8694 505494
rect -8458 505258 -8374 505494
rect -8138 505258 -8106 505494
rect -8726 505174 -8106 505258
rect -8726 504938 -8694 505174
rect -8458 504938 -8374 505174
rect -8138 504938 -8106 505174
rect -8726 471494 -8106 504938
rect -8726 471258 -8694 471494
rect -8458 471258 -8374 471494
rect -8138 471258 -8106 471494
rect -8726 471174 -8106 471258
rect -8726 470938 -8694 471174
rect -8458 470938 -8374 471174
rect -8138 470938 -8106 471174
rect -8726 437494 -8106 470938
rect -8726 437258 -8694 437494
rect -8458 437258 -8374 437494
rect -8138 437258 -8106 437494
rect -8726 437174 -8106 437258
rect -8726 436938 -8694 437174
rect -8458 436938 -8374 437174
rect -8138 436938 -8106 437174
rect -8726 403494 -8106 436938
rect -8726 403258 -8694 403494
rect -8458 403258 -8374 403494
rect -8138 403258 -8106 403494
rect -8726 403174 -8106 403258
rect -8726 402938 -8694 403174
rect -8458 402938 -8374 403174
rect -8138 402938 -8106 403174
rect -8726 369494 -8106 402938
rect -8726 369258 -8694 369494
rect -8458 369258 -8374 369494
rect -8138 369258 -8106 369494
rect -8726 369174 -8106 369258
rect -8726 368938 -8694 369174
rect -8458 368938 -8374 369174
rect -8138 368938 -8106 369174
rect -8726 335494 -8106 368938
rect -8726 335258 -8694 335494
rect -8458 335258 -8374 335494
rect -8138 335258 -8106 335494
rect -8726 335174 -8106 335258
rect -8726 334938 -8694 335174
rect -8458 334938 -8374 335174
rect -8138 334938 -8106 335174
rect -8726 301494 -8106 334938
rect -8726 301258 -8694 301494
rect -8458 301258 -8374 301494
rect -8138 301258 -8106 301494
rect -8726 301174 -8106 301258
rect -8726 300938 -8694 301174
rect -8458 300938 -8374 301174
rect -8138 300938 -8106 301174
rect -8726 267494 -8106 300938
rect -8726 267258 -8694 267494
rect -8458 267258 -8374 267494
rect -8138 267258 -8106 267494
rect -8726 267174 -8106 267258
rect -8726 266938 -8694 267174
rect -8458 266938 -8374 267174
rect -8138 266938 -8106 267174
rect -8726 233494 -8106 266938
rect -8726 233258 -8694 233494
rect -8458 233258 -8374 233494
rect -8138 233258 -8106 233494
rect -8726 233174 -8106 233258
rect -8726 232938 -8694 233174
rect -8458 232938 -8374 233174
rect -8138 232938 -8106 233174
rect -8726 199494 -8106 232938
rect -8726 199258 -8694 199494
rect -8458 199258 -8374 199494
rect -8138 199258 -8106 199494
rect -8726 199174 -8106 199258
rect -8726 198938 -8694 199174
rect -8458 198938 -8374 199174
rect -8138 198938 -8106 199174
rect -8726 165494 -8106 198938
rect -8726 165258 -8694 165494
rect -8458 165258 -8374 165494
rect -8138 165258 -8106 165494
rect -8726 165174 -8106 165258
rect -8726 164938 -8694 165174
rect -8458 164938 -8374 165174
rect -8138 164938 -8106 165174
rect -8726 131494 -8106 164938
rect -8726 131258 -8694 131494
rect -8458 131258 -8374 131494
rect -8138 131258 -8106 131494
rect -8726 131174 -8106 131258
rect -8726 130938 -8694 131174
rect -8458 130938 -8374 131174
rect -8138 130938 -8106 131174
rect -8726 97494 -8106 130938
rect -8726 97258 -8694 97494
rect -8458 97258 -8374 97494
rect -8138 97258 -8106 97494
rect -8726 97174 -8106 97258
rect -8726 96938 -8694 97174
rect -8458 96938 -8374 97174
rect -8138 96938 -8106 97174
rect -8726 63494 -8106 96938
rect -8726 63258 -8694 63494
rect -8458 63258 -8374 63494
rect -8138 63258 -8106 63494
rect -8726 63174 -8106 63258
rect -8726 62938 -8694 63174
rect -8458 62938 -8374 63174
rect -8138 62938 -8106 63174
rect -8726 29494 -8106 62938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 671774 -7146 710042
rect -7766 671538 -7734 671774
rect -7498 671538 -7414 671774
rect -7178 671538 -7146 671774
rect -7766 671454 -7146 671538
rect -7766 671218 -7734 671454
rect -7498 671218 -7414 671454
rect -7178 671218 -7146 671454
rect -7766 637774 -7146 671218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 603774 -7146 637218
rect -7766 603538 -7734 603774
rect -7498 603538 -7414 603774
rect -7178 603538 -7146 603774
rect -7766 603454 -7146 603538
rect -7766 603218 -7734 603454
rect -7498 603218 -7414 603454
rect -7178 603218 -7146 603454
rect -7766 569774 -7146 603218
rect -7766 569538 -7734 569774
rect -7498 569538 -7414 569774
rect -7178 569538 -7146 569774
rect -7766 569454 -7146 569538
rect -7766 569218 -7734 569454
rect -7498 569218 -7414 569454
rect -7178 569218 -7146 569454
rect -7766 535774 -7146 569218
rect -7766 535538 -7734 535774
rect -7498 535538 -7414 535774
rect -7178 535538 -7146 535774
rect -7766 535454 -7146 535538
rect -7766 535218 -7734 535454
rect -7498 535218 -7414 535454
rect -7178 535218 -7146 535454
rect -7766 501774 -7146 535218
rect -7766 501538 -7734 501774
rect -7498 501538 -7414 501774
rect -7178 501538 -7146 501774
rect -7766 501454 -7146 501538
rect -7766 501218 -7734 501454
rect -7498 501218 -7414 501454
rect -7178 501218 -7146 501454
rect -7766 467774 -7146 501218
rect -7766 467538 -7734 467774
rect -7498 467538 -7414 467774
rect -7178 467538 -7146 467774
rect -7766 467454 -7146 467538
rect -7766 467218 -7734 467454
rect -7498 467218 -7414 467454
rect -7178 467218 -7146 467454
rect -7766 433774 -7146 467218
rect -7766 433538 -7734 433774
rect -7498 433538 -7414 433774
rect -7178 433538 -7146 433774
rect -7766 433454 -7146 433538
rect -7766 433218 -7734 433454
rect -7498 433218 -7414 433454
rect -7178 433218 -7146 433454
rect -7766 399774 -7146 433218
rect -7766 399538 -7734 399774
rect -7498 399538 -7414 399774
rect -7178 399538 -7146 399774
rect -7766 399454 -7146 399538
rect -7766 399218 -7734 399454
rect -7498 399218 -7414 399454
rect -7178 399218 -7146 399454
rect -7766 365774 -7146 399218
rect -7766 365538 -7734 365774
rect -7498 365538 -7414 365774
rect -7178 365538 -7146 365774
rect -7766 365454 -7146 365538
rect -7766 365218 -7734 365454
rect -7498 365218 -7414 365454
rect -7178 365218 -7146 365454
rect -7766 331774 -7146 365218
rect -7766 331538 -7734 331774
rect -7498 331538 -7414 331774
rect -7178 331538 -7146 331774
rect -7766 331454 -7146 331538
rect -7766 331218 -7734 331454
rect -7498 331218 -7414 331454
rect -7178 331218 -7146 331454
rect -7766 297774 -7146 331218
rect -7766 297538 -7734 297774
rect -7498 297538 -7414 297774
rect -7178 297538 -7146 297774
rect -7766 297454 -7146 297538
rect -7766 297218 -7734 297454
rect -7498 297218 -7414 297454
rect -7178 297218 -7146 297454
rect -7766 263774 -7146 297218
rect -7766 263538 -7734 263774
rect -7498 263538 -7414 263774
rect -7178 263538 -7146 263774
rect -7766 263454 -7146 263538
rect -7766 263218 -7734 263454
rect -7498 263218 -7414 263454
rect -7178 263218 -7146 263454
rect -7766 229774 -7146 263218
rect -7766 229538 -7734 229774
rect -7498 229538 -7414 229774
rect -7178 229538 -7146 229774
rect -7766 229454 -7146 229538
rect -7766 229218 -7734 229454
rect -7498 229218 -7414 229454
rect -7178 229218 -7146 229454
rect -7766 195774 -7146 229218
rect -7766 195538 -7734 195774
rect -7498 195538 -7414 195774
rect -7178 195538 -7146 195774
rect -7766 195454 -7146 195538
rect -7766 195218 -7734 195454
rect -7498 195218 -7414 195454
rect -7178 195218 -7146 195454
rect -7766 161774 -7146 195218
rect -7766 161538 -7734 161774
rect -7498 161538 -7414 161774
rect -7178 161538 -7146 161774
rect -7766 161454 -7146 161538
rect -7766 161218 -7734 161454
rect -7498 161218 -7414 161454
rect -7178 161218 -7146 161454
rect -7766 127774 -7146 161218
rect -7766 127538 -7734 127774
rect -7498 127538 -7414 127774
rect -7178 127538 -7146 127774
rect -7766 127454 -7146 127538
rect -7766 127218 -7734 127454
rect -7498 127218 -7414 127454
rect -7178 127218 -7146 127454
rect -7766 93774 -7146 127218
rect -7766 93538 -7734 93774
rect -7498 93538 -7414 93774
rect -7178 93538 -7146 93774
rect -7766 93454 -7146 93538
rect -7766 93218 -7734 93454
rect -7498 93218 -7414 93454
rect -7178 93218 -7146 93454
rect -7766 59774 -7146 93218
rect -7766 59538 -7734 59774
rect -7498 59538 -7414 59774
rect -7178 59538 -7146 59774
rect -7766 59454 -7146 59538
rect -7766 59218 -7734 59454
rect -7498 59218 -7414 59454
rect -7178 59218 -7146 59454
rect -7766 25774 -7146 59218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 668054 -6186 709082
rect -6806 667818 -6774 668054
rect -6538 667818 -6454 668054
rect -6218 667818 -6186 668054
rect -6806 667734 -6186 667818
rect -6806 667498 -6774 667734
rect -6538 667498 -6454 667734
rect -6218 667498 -6186 667734
rect -6806 634054 -6186 667498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 600054 -6186 633498
rect -6806 599818 -6774 600054
rect -6538 599818 -6454 600054
rect -6218 599818 -6186 600054
rect -6806 599734 -6186 599818
rect -6806 599498 -6774 599734
rect -6538 599498 -6454 599734
rect -6218 599498 -6186 599734
rect -6806 566054 -6186 599498
rect -6806 565818 -6774 566054
rect -6538 565818 -6454 566054
rect -6218 565818 -6186 566054
rect -6806 565734 -6186 565818
rect -6806 565498 -6774 565734
rect -6538 565498 -6454 565734
rect -6218 565498 -6186 565734
rect -6806 532054 -6186 565498
rect -6806 531818 -6774 532054
rect -6538 531818 -6454 532054
rect -6218 531818 -6186 532054
rect -6806 531734 -6186 531818
rect -6806 531498 -6774 531734
rect -6538 531498 -6454 531734
rect -6218 531498 -6186 531734
rect -6806 498054 -6186 531498
rect -6806 497818 -6774 498054
rect -6538 497818 -6454 498054
rect -6218 497818 -6186 498054
rect -6806 497734 -6186 497818
rect -6806 497498 -6774 497734
rect -6538 497498 -6454 497734
rect -6218 497498 -6186 497734
rect -6806 464054 -6186 497498
rect -6806 463818 -6774 464054
rect -6538 463818 -6454 464054
rect -6218 463818 -6186 464054
rect -6806 463734 -6186 463818
rect -6806 463498 -6774 463734
rect -6538 463498 -6454 463734
rect -6218 463498 -6186 463734
rect -6806 430054 -6186 463498
rect -6806 429818 -6774 430054
rect -6538 429818 -6454 430054
rect -6218 429818 -6186 430054
rect -6806 429734 -6186 429818
rect -6806 429498 -6774 429734
rect -6538 429498 -6454 429734
rect -6218 429498 -6186 429734
rect -6806 396054 -6186 429498
rect -6806 395818 -6774 396054
rect -6538 395818 -6454 396054
rect -6218 395818 -6186 396054
rect -6806 395734 -6186 395818
rect -6806 395498 -6774 395734
rect -6538 395498 -6454 395734
rect -6218 395498 -6186 395734
rect -6806 362054 -6186 395498
rect -6806 361818 -6774 362054
rect -6538 361818 -6454 362054
rect -6218 361818 -6186 362054
rect -6806 361734 -6186 361818
rect -6806 361498 -6774 361734
rect -6538 361498 -6454 361734
rect -6218 361498 -6186 361734
rect -6806 328054 -6186 361498
rect -6806 327818 -6774 328054
rect -6538 327818 -6454 328054
rect -6218 327818 -6186 328054
rect -6806 327734 -6186 327818
rect -6806 327498 -6774 327734
rect -6538 327498 -6454 327734
rect -6218 327498 -6186 327734
rect -6806 294054 -6186 327498
rect -6806 293818 -6774 294054
rect -6538 293818 -6454 294054
rect -6218 293818 -6186 294054
rect -6806 293734 -6186 293818
rect -6806 293498 -6774 293734
rect -6538 293498 -6454 293734
rect -6218 293498 -6186 293734
rect -6806 260054 -6186 293498
rect -6806 259818 -6774 260054
rect -6538 259818 -6454 260054
rect -6218 259818 -6186 260054
rect -6806 259734 -6186 259818
rect -6806 259498 -6774 259734
rect -6538 259498 -6454 259734
rect -6218 259498 -6186 259734
rect -6806 226054 -6186 259498
rect -6806 225818 -6774 226054
rect -6538 225818 -6454 226054
rect -6218 225818 -6186 226054
rect -6806 225734 -6186 225818
rect -6806 225498 -6774 225734
rect -6538 225498 -6454 225734
rect -6218 225498 -6186 225734
rect -6806 192054 -6186 225498
rect -6806 191818 -6774 192054
rect -6538 191818 -6454 192054
rect -6218 191818 -6186 192054
rect -6806 191734 -6186 191818
rect -6806 191498 -6774 191734
rect -6538 191498 -6454 191734
rect -6218 191498 -6186 191734
rect -6806 158054 -6186 191498
rect -6806 157818 -6774 158054
rect -6538 157818 -6454 158054
rect -6218 157818 -6186 158054
rect -6806 157734 -6186 157818
rect -6806 157498 -6774 157734
rect -6538 157498 -6454 157734
rect -6218 157498 -6186 157734
rect -6806 124054 -6186 157498
rect -6806 123818 -6774 124054
rect -6538 123818 -6454 124054
rect -6218 123818 -6186 124054
rect -6806 123734 -6186 123818
rect -6806 123498 -6774 123734
rect -6538 123498 -6454 123734
rect -6218 123498 -6186 123734
rect -6806 90054 -6186 123498
rect -6806 89818 -6774 90054
rect -6538 89818 -6454 90054
rect -6218 89818 -6186 90054
rect -6806 89734 -6186 89818
rect -6806 89498 -6774 89734
rect -6538 89498 -6454 89734
rect -6218 89498 -6186 89734
rect -6806 56054 -6186 89498
rect -6806 55818 -6774 56054
rect -6538 55818 -6454 56054
rect -6218 55818 -6186 56054
rect -6806 55734 -6186 55818
rect -6806 55498 -6774 55734
rect -6538 55498 -6454 55734
rect -6218 55498 -6186 55734
rect -6806 22054 -6186 55498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 698334 -5226 708122
rect -5846 698098 -5814 698334
rect -5578 698098 -5494 698334
rect -5258 698098 -5226 698334
rect -5846 698014 -5226 698098
rect -5846 697778 -5814 698014
rect -5578 697778 -5494 698014
rect -5258 697778 -5226 698014
rect -5846 664334 -5226 697778
rect -5846 664098 -5814 664334
rect -5578 664098 -5494 664334
rect -5258 664098 -5226 664334
rect -5846 664014 -5226 664098
rect -5846 663778 -5814 664014
rect -5578 663778 -5494 664014
rect -5258 663778 -5226 664014
rect -5846 630334 -5226 663778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 596334 -5226 629778
rect -5846 596098 -5814 596334
rect -5578 596098 -5494 596334
rect -5258 596098 -5226 596334
rect -5846 596014 -5226 596098
rect -5846 595778 -5814 596014
rect -5578 595778 -5494 596014
rect -5258 595778 -5226 596014
rect -5846 562334 -5226 595778
rect -5846 562098 -5814 562334
rect -5578 562098 -5494 562334
rect -5258 562098 -5226 562334
rect -5846 562014 -5226 562098
rect -5846 561778 -5814 562014
rect -5578 561778 -5494 562014
rect -5258 561778 -5226 562014
rect -5846 528334 -5226 561778
rect -5846 528098 -5814 528334
rect -5578 528098 -5494 528334
rect -5258 528098 -5226 528334
rect -5846 528014 -5226 528098
rect -5846 527778 -5814 528014
rect -5578 527778 -5494 528014
rect -5258 527778 -5226 528014
rect -5846 494334 -5226 527778
rect -5846 494098 -5814 494334
rect -5578 494098 -5494 494334
rect -5258 494098 -5226 494334
rect -5846 494014 -5226 494098
rect -5846 493778 -5814 494014
rect -5578 493778 -5494 494014
rect -5258 493778 -5226 494014
rect -5846 460334 -5226 493778
rect -5846 460098 -5814 460334
rect -5578 460098 -5494 460334
rect -5258 460098 -5226 460334
rect -5846 460014 -5226 460098
rect -5846 459778 -5814 460014
rect -5578 459778 -5494 460014
rect -5258 459778 -5226 460014
rect -5846 426334 -5226 459778
rect -5846 426098 -5814 426334
rect -5578 426098 -5494 426334
rect -5258 426098 -5226 426334
rect -5846 426014 -5226 426098
rect -5846 425778 -5814 426014
rect -5578 425778 -5494 426014
rect -5258 425778 -5226 426014
rect -5846 392334 -5226 425778
rect -5846 392098 -5814 392334
rect -5578 392098 -5494 392334
rect -5258 392098 -5226 392334
rect -5846 392014 -5226 392098
rect -5846 391778 -5814 392014
rect -5578 391778 -5494 392014
rect -5258 391778 -5226 392014
rect -5846 358334 -5226 391778
rect -5846 358098 -5814 358334
rect -5578 358098 -5494 358334
rect -5258 358098 -5226 358334
rect -5846 358014 -5226 358098
rect -5846 357778 -5814 358014
rect -5578 357778 -5494 358014
rect -5258 357778 -5226 358014
rect -5846 324334 -5226 357778
rect -5846 324098 -5814 324334
rect -5578 324098 -5494 324334
rect -5258 324098 -5226 324334
rect -5846 324014 -5226 324098
rect -5846 323778 -5814 324014
rect -5578 323778 -5494 324014
rect -5258 323778 -5226 324014
rect -5846 290334 -5226 323778
rect -5846 290098 -5814 290334
rect -5578 290098 -5494 290334
rect -5258 290098 -5226 290334
rect -5846 290014 -5226 290098
rect -5846 289778 -5814 290014
rect -5578 289778 -5494 290014
rect -5258 289778 -5226 290014
rect -5846 256334 -5226 289778
rect -5846 256098 -5814 256334
rect -5578 256098 -5494 256334
rect -5258 256098 -5226 256334
rect -5846 256014 -5226 256098
rect -5846 255778 -5814 256014
rect -5578 255778 -5494 256014
rect -5258 255778 -5226 256014
rect -5846 222334 -5226 255778
rect -5846 222098 -5814 222334
rect -5578 222098 -5494 222334
rect -5258 222098 -5226 222334
rect -5846 222014 -5226 222098
rect -5846 221778 -5814 222014
rect -5578 221778 -5494 222014
rect -5258 221778 -5226 222014
rect -5846 188334 -5226 221778
rect -5846 188098 -5814 188334
rect -5578 188098 -5494 188334
rect -5258 188098 -5226 188334
rect -5846 188014 -5226 188098
rect -5846 187778 -5814 188014
rect -5578 187778 -5494 188014
rect -5258 187778 -5226 188014
rect -5846 154334 -5226 187778
rect -5846 154098 -5814 154334
rect -5578 154098 -5494 154334
rect -5258 154098 -5226 154334
rect -5846 154014 -5226 154098
rect -5846 153778 -5814 154014
rect -5578 153778 -5494 154014
rect -5258 153778 -5226 154014
rect -5846 120334 -5226 153778
rect -5846 120098 -5814 120334
rect -5578 120098 -5494 120334
rect -5258 120098 -5226 120334
rect -5846 120014 -5226 120098
rect -5846 119778 -5814 120014
rect -5578 119778 -5494 120014
rect -5258 119778 -5226 120014
rect -5846 86334 -5226 119778
rect -5846 86098 -5814 86334
rect -5578 86098 -5494 86334
rect -5258 86098 -5226 86334
rect -5846 86014 -5226 86098
rect -5846 85778 -5814 86014
rect -5578 85778 -5494 86014
rect -5258 85778 -5226 86014
rect -5846 52334 -5226 85778
rect -5846 52098 -5814 52334
rect -5578 52098 -5494 52334
rect -5258 52098 -5226 52334
rect -5846 52014 -5226 52098
rect -5846 51778 -5814 52014
rect -5578 51778 -5494 52014
rect -5258 51778 -5226 52014
rect -5846 18334 -5226 51778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 694614 -4266 707162
rect -4886 694378 -4854 694614
rect -4618 694378 -4534 694614
rect -4298 694378 -4266 694614
rect -4886 694294 -4266 694378
rect -4886 694058 -4854 694294
rect -4618 694058 -4534 694294
rect -4298 694058 -4266 694294
rect -4886 660614 -4266 694058
rect -4886 660378 -4854 660614
rect -4618 660378 -4534 660614
rect -4298 660378 -4266 660614
rect -4886 660294 -4266 660378
rect -4886 660058 -4854 660294
rect -4618 660058 -4534 660294
rect -4298 660058 -4266 660294
rect -4886 626614 -4266 660058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 592614 -4266 626058
rect -4886 592378 -4854 592614
rect -4618 592378 -4534 592614
rect -4298 592378 -4266 592614
rect -4886 592294 -4266 592378
rect -4886 592058 -4854 592294
rect -4618 592058 -4534 592294
rect -4298 592058 -4266 592294
rect -4886 558614 -4266 592058
rect -4886 558378 -4854 558614
rect -4618 558378 -4534 558614
rect -4298 558378 -4266 558614
rect -4886 558294 -4266 558378
rect -4886 558058 -4854 558294
rect -4618 558058 -4534 558294
rect -4298 558058 -4266 558294
rect -4886 524614 -4266 558058
rect -4886 524378 -4854 524614
rect -4618 524378 -4534 524614
rect -4298 524378 -4266 524614
rect -4886 524294 -4266 524378
rect -4886 524058 -4854 524294
rect -4618 524058 -4534 524294
rect -4298 524058 -4266 524294
rect -4886 490614 -4266 524058
rect -4886 490378 -4854 490614
rect -4618 490378 -4534 490614
rect -4298 490378 -4266 490614
rect -4886 490294 -4266 490378
rect -4886 490058 -4854 490294
rect -4618 490058 -4534 490294
rect -4298 490058 -4266 490294
rect -4886 456614 -4266 490058
rect -4886 456378 -4854 456614
rect -4618 456378 -4534 456614
rect -4298 456378 -4266 456614
rect -4886 456294 -4266 456378
rect -4886 456058 -4854 456294
rect -4618 456058 -4534 456294
rect -4298 456058 -4266 456294
rect -4886 422614 -4266 456058
rect -4886 422378 -4854 422614
rect -4618 422378 -4534 422614
rect -4298 422378 -4266 422614
rect -4886 422294 -4266 422378
rect -4886 422058 -4854 422294
rect -4618 422058 -4534 422294
rect -4298 422058 -4266 422294
rect -4886 388614 -4266 422058
rect -4886 388378 -4854 388614
rect -4618 388378 -4534 388614
rect -4298 388378 -4266 388614
rect -4886 388294 -4266 388378
rect -4886 388058 -4854 388294
rect -4618 388058 -4534 388294
rect -4298 388058 -4266 388294
rect -4886 354614 -4266 388058
rect -4886 354378 -4854 354614
rect -4618 354378 -4534 354614
rect -4298 354378 -4266 354614
rect -4886 354294 -4266 354378
rect -4886 354058 -4854 354294
rect -4618 354058 -4534 354294
rect -4298 354058 -4266 354294
rect -4886 320614 -4266 354058
rect -4886 320378 -4854 320614
rect -4618 320378 -4534 320614
rect -4298 320378 -4266 320614
rect -4886 320294 -4266 320378
rect -4886 320058 -4854 320294
rect -4618 320058 -4534 320294
rect -4298 320058 -4266 320294
rect -4886 286614 -4266 320058
rect -4886 286378 -4854 286614
rect -4618 286378 -4534 286614
rect -4298 286378 -4266 286614
rect -4886 286294 -4266 286378
rect -4886 286058 -4854 286294
rect -4618 286058 -4534 286294
rect -4298 286058 -4266 286294
rect -4886 252614 -4266 286058
rect -4886 252378 -4854 252614
rect -4618 252378 -4534 252614
rect -4298 252378 -4266 252614
rect -4886 252294 -4266 252378
rect -4886 252058 -4854 252294
rect -4618 252058 -4534 252294
rect -4298 252058 -4266 252294
rect -4886 218614 -4266 252058
rect -4886 218378 -4854 218614
rect -4618 218378 -4534 218614
rect -4298 218378 -4266 218614
rect -4886 218294 -4266 218378
rect -4886 218058 -4854 218294
rect -4618 218058 -4534 218294
rect -4298 218058 -4266 218294
rect -4886 184614 -4266 218058
rect -4886 184378 -4854 184614
rect -4618 184378 -4534 184614
rect -4298 184378 -4266 184614
rect -4886 184294 -4266 184378
rect -4886 184058 -4854 184294
rect -4618 184058 -4534 184294
rect -4298 184058 -4266 184294
rect -4886 150614 -4266 184058
rect -4886 150378 -4854 150614
rect -4618 150378 -4534 150614
rect -4298 150378 -4266 150614
rect -4886 150294 -4266 150378
rect -4886 150058 -4854 150294
rect -4618 150058 -4534 150294
rect -4298 150058 -4266 150294
rect -4886 116614 -4266 150058
rect -4886 116378 -4854 116614
rect -4618 116378 -4534 116614
rect -4298 116378 -4266 116614
rect -4886 116294 -4266 116378
rect -4886 116058 -4854 116294
rect -4618 116058 -4534 116294
rect -4298 116058 -4266 116294
rect -4886 82614 -4266 116058
rect -4886 82378 -4854 82614
rect -4618 82378 -4534 82614
rect -4298 82378 -4266 82614
rect -4886 82294 -4266 82378
rect -4886 82058 -4854 82294
rect -4618 82058 -4534 82294
rect -4298 82058 -4266 82294
rect -4886 48614 -4266 82058
rect -4886 48378 -4854 48614
rect -4618 48378 -4534 48614
rect -4298 48378 -4266 48614
rect -4886 48294 -4266 48378
rect -4886 48058 -4854 48294
rect -4618 48058 -4534 48294
rect -4298 48058 -4266 48294
rect -4886 14614 -4266 48058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 690894 -3306 706202
rect -3926 690658 -3894 690894
rect -3658 690658 -3574 690894
rect -3338 690658 -3306 690894
rect -3926 690574 -3306 690658
rect -3926 690338 -3894 690574
rect -3658 690338 -3574 690574
rect -3338 690338 -3306 690574
rect -3926 656894 -3306 690338
rect -3926 656658 -3894 656894
rect -3658 656658 -3574 656894
rect -3338 656658 -3306 656894
rect -3926 656574 -3306 656658
rect -3926 656338 -3894 656574
rect -3658 656338 -3574 656574
rect -3338 656338 -3306 656574
rect -3926 622894 -3306 656338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 588894 -3306 622338
rect -3926 588658 -3894 588894
rect -3658 588658 -3574 588894
rect -3338 588658 -3306 588894
rect -3926 588574 -3306 588658
rect -3926 588338 -3894 588574
rect -3658 588338 -3574 588574
rect -3338 588338 -3306 588574
rect -3926 554894 -3306 588338
rect -3926 554658 -3894 554894
rect -3658 554658 -3574 554894
rect -3338 554658 -3306 554894
rect -3926 554574 -3306 554658
rect -3926 554338 -3894 554574
rect -3658 554338 -3574 554574
rect -3338 554338 -3306 554574
rect -3926 520894 -3306 554338
rect -3926 520658 -3894 520894
rect -3658 520658 -3574 520894
rect -3338 520658 -3306 520894
rect -3926 520574 -3306 520658
rect -3926 520338 -3894 520574
rect -3658 520338 -3574 520574
rect -3338 520338 -3306 520574
rect -3926 486894 -3306 520338
rect -3926 486658 -3894 486894
rect -3658 486658 -3574 486894
rect -3338 486658 -3306 486894
rect -3926 486574 -3306 486658
rect -3926 486338 -3894 486574
rect -3658 486338 -3574 486574
rect -3338 486338 -3306 486574
rect -3926 452894 -3306 486338
rect -3926 452658 -3894 452894
rect -3658 452658 -3574 452894
rect -3338 452658 -3306 452894
rect -3926 452574 -3306 452658
rect -3926 452338 -3894 452574
rect -3658 452338 -3574 452574
rect -3338 452338 -3306 452574
rect -3926 418894 -3306 452338
rect -3926 418658 -3894 418894
rect -3658 418658 -3574 418894
rect -3338 418658 -3306 418894
rect -3926 418574 -3306 418658
rect -3926 418338 -3894 418574
rect -3658 418338 -3574 418574
rect -3338 418338 -3306 418574
rect -3926 384894 -3306 418338
rect -3926 384658 -3894 384894
rect -3658 384658 -3574 384894
rect -3338 384658 -3306 384894
rect -3926 384574 -3306 384658
rect -3926 384338 -3894 384574
rect -3658 384338 -3574 384574
rect -3338 384338 -3306 384574
rect -3926 350894 -3306 384338
rect -3926 350658 -3894 350894
rect -3658 350658 -3574 350894
rect -3338 350658 -3306 350894
rect -3926 350574 -3306 350658
rect -3926 350338 -3894 350574
rect -3658 350338 -3574 350574
rect -3338 350338 -3306 350574
rect -3926 316894 -3306 350338
rect -3926 316658 -3894 316894
rect -3658 316658 -3574 316894
rect -3338 316658 -3306 316894
rect -3926 316574 -3306 316658
rect -3926 316338 -3894 316574
rect -3658 316338 -3574 316574
rect -3338 316338 -3306 316574
rect -3926 282894 -3306 316338
rect -3926 282658 -3894 282894
rect -3658 282658 -3574 282894
rect -3338 282658 -3306 282894
rect -3926 282574 -3306 282658
rect -3926 282338 -3894 282574
rect -3658 282338 -3574 282574
rect -3338 282338 -3306 282574
rect -3926 248894 -3306 282338
rect -3926 248658 -3894 248894
rect -3658 248658 -3574 248894
rect -3338 248658 -3306 248894
rect -3926 248574 -3306 248658
rect -3926 248338 -3894 248574
rect -3658 248338 -3574 248574
rect -3338 248338 -3306 248574
rect -3926 214894 -3306 248338
rect -3926 214658 -3894 214894
rect -3658 214658 -3574 214894
rect -3338 214658 -3306 214894
rect -3926 214574 -3306 214658
rect -3926 214338 -3894 214574
rect -3658 214338 -3574 214574
rect -3338 214338 -3306 214574
rect -3926 180894 -3306 214338
rect -3926 180658 -3894 180894
rect -3658 180658 -3574 180894
rect -3338 180658 -3306 180894
rect -3926 180574 -3306 180658
rect -3926 180338 -3894 180574
rect -3658 180338 -3574 180574
rect -3338 180338 -3306 180574
rect -3926 146894 -3306 180338
rect -3926 146658 -3894 146894
rect -3658 146658 -3574 146894
rect -3338 146658 -3306 146894
rect -3926 146574 -3306 146658
rect -3926 146338 -3894 146574
rect -3658 146338 -3574 146574
rect -3338 146338 -3306 146574
rect -3926 112894 -3306 146338
rect -3926 112658 -3894 112894
rect -3658 112658 -3574 112894
rect -3338 112658 -3306 112894
rect -3926 112574 -3306 112658
rect -3926 112338 -3894 112574
rect -3658 112338 -3574 112574
rect -3338 112338 -3306 112574
rect -3926 78894 -3306 112338
rect -3926 78658 -3894 78894
rect -3658 78658 -3574 78894
rect -3338 78658 -3306 78894
rect -3926 78574 -3306 78658
rect -3926 78338 -3894 78574
rect -3658 78338 -3574 78574
rect -3338 78338 -3306 78574
rect -3926 44894 -3306 78338
rect -3926 44658 -3894 44894
rect -3658 44658 -3574 44894
rect -3338 44658 -3306 44894
rect -3926 44574 -3306 44658
rect -3926 44338 -3894 44574
rect -3658 44338 -3574 44574
rect -3338 44338 -3306 44574
rect -3926 10894 -3306 44338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 687174 -2346 705242
rect -2966 686938 -2934 687174
rect -2698 686938 -2614 687174
rect -2378 686938 -2346 687174
rect -2966 686854 -2346 686938
rect -2966 686618 -2934 686854
rect -2698 686618 -2614 686854
rect -2378 686618 -2346 686854
rect -2966 653174 -2346 686618
rect -2966 652938 -2934 653174
rect -2698 652938 -2614 653174
rect -2378 652938 -2346 653174
rect -2966 652854 -2346 652938
rect -2966 652618 -2934 652854
rect -2698 652618 -2614 652854
rect -2378 652618 -2346 652854
rect -2966 619174 -2346 652618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 585174 -2346 618618
rect -2966 584938 -2934 585174
rect -2698 584938 -2614 585174
rect -2378 584938 -2346 585174
rect -2966 584854 -2346 584938
rect -2966 584618 -2934 584854
rect -2698 584618 -2614 584854
rect -2378 584618 -2346 584854
rect -2966 551174 -2346 584618
rect -2966 550938 -2934 551174
rect -2698 550938 -2614 551174
rect -2378 550938 -2346 551174
rect -2966 550854 -2346 550938
rect -2966 550618 -2934 550854
rect -2698 550618 -2614 550854
rect -2378 550618 -2346 550854
rect -2966 517174 -2346 550618
rect -2966 516938 -2934 517174
rect -2698 516938 -2614 517174
rect -2378 516938 -2346 517174
rect -2966 516854 -2346 516938
rect -2966 516618 -2934 516854
rect -2698 516618 -2614 516854
rect -2378 516618 -2346 516854
rect -2966 483174 -2346 516618
rect -2966 482938 -2934 483174
rect -2698 482938 -2614 483174
rect -2378 482938 -2346 483174
rect -2966 482854 -2346 482938
rect -2966 482618 -2934 482854
rect -2698 482618 -2614 482854
rect -2378 482618 -2346 482854
rect -2966 449174 -2346 482618
rect -2966 448938 -2934 449174
rect -2698 448938 -2614 449174
rect -2378 448938 -2346 449174
rect -2966 448854 -2346 448938
rect -2966 448618 -2934 448854
rect -2698 448618 -2614 448854
rect -2378 448618 -2346 448854
rect -2966 415174 -2346 448618
rect -2966 414938 -2934 415174
rect -2698 414938 -2614 415174
rect -2378 414938 -2346 415174
rect -2966 414854 -2346 414938
rect -2966 414618 -2934 414854
rect -2698 414618 -2614 414854
rect -2378 414618 -2346 414854
rect -2966 381174 -2346 414618
rect -2966 380938 -2934 381174
rect -2698 380938 -2614 381174
rect -2378 380938 -2346 381174
rect -2966 380854 -2346 380938
rect -2966 380618 -2934 380854
rect -2698 380618 -2614 380854
rect -2378 380618 -2346 380854
rect -2966 347174 -2346 380618
rect -2966 346938 -2934 347174
rect -2698 346938 -2614 347174
rect -2378 346938 -2346 347174
rect -2966 346854 -2346 346938
rect -2966 346618 -2934 346854
rect -2698 346618 -2614 346854
rect -2378 346618 -2346 346854
rect -2966 313174 -2346 346618
rect -2966 312938 -2934 313174
rect -2698 312938 -2614 313174
rect -2378 312938 -2346 313174
rect -2966 312854 -2346 312938
rect -2966 312618 -2934 312854
rect -2698 312618 -2614 312854
rect -2378 312618 -2346 312854
rect -2966 279174 -2346 312618
rect -2966 278938 -2934 279174
rect -2698 278938 -2614 279174
rect -2378 278938 -2346 279174
rect -2966 278854 -2346 278938
rect -2966 278618 -2934 278854
rect -2698 278618 -2614 278854
rect -2378 278618 -2346 278854
rect -2966 245174 -2346 278618
rect -2966 244938 -2934 245174
rect -2698 244938 -2614 245174
rect -2378 244938 -2346 245174
rect -2966 244854 -2346 244938
rect -2966 244618 -2934 244854
rect -2698 244618 -2614 244854
rect -2378 244618 -2346 244854
rect -2966 211174 -2346 244618
rect -2966 210938 -2934 211174
rect -2698 210938 -2614 211174
rect -2378 210938 -2346 211174
rect -2966 210854 -2346 210938
rect -2966 210618 -2934 210854
rect -2698 210618 -2614 210854
rect -2378 210618 -2346 210854
rect -2966 177174 -2346 210618
rect -2966 176938 -2934 177174
rect -2698 176938 -2614 177174
rect -2378 176938 -2346 177174
rect -2966 176854 -2346 176938
rect -2966 176618 -2934 176854
rect -2698 176618 -2614 176854
rect -2378 176618 -2346 176854
rect -2966 143174 -2346 176618
rect -2966 142938 -2934 143174
rect -2698 142938 -2614 143174
rect -2378 142938 -2346 143174
rect -2966 142854 -2346 142938
rect -2966 142618 -2934 142854
rect -2698 142618 -2614 142854
rect -2378 142618 -2346 142854
rect -2966 109174 -2346 142618
rect -2966 108938 -2934 109174
rect -2698 108938 -2614 109174
rect -2378 108938 -2346 109174
rect -2966 108854 -2346 108938
rect -2966 108618 -2934 108854
rect -2698 108618 -2614 108854
rect -2378 108618 -2346 108854
rect -2966 75174 -2346 108618
rect -2966 74938 -2934 75174
rect -2698 74938 -2614 75174
rect -2378 74938 -2346 75174
rect -2966 74854 -2346 74938
rect -2966 74618 -2934 74854
rect -2698 74618 -2614 74854
rect -2378 74618 -2346 74854
rect -2966 41174 -2346 74618
rect -2966 40938 -2934 41174
rect -2698 40938 -2614 41174
rect -2378 40938 -2346 41174
rect -2966 40854 -2346 40938
rect -2966 40618 -2934 40854
rect -2698 40618 -2614 40854
rect -2378 40618 -2346 40854
rect -2966 7174 -2346 40618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 683454 -1386 704282
rect -2006 683218 -1974 683454
rect -1738 683218 -1654 683454
rect -1418 683218 -1386 683454
rect -2006 683134 -1386 683218
rect -2006 682898 -1974 683134
rect -1738 682898 -1654 683134
rect -1418 682898 -1386 683134
rect -2006 649454 -1386 682898
rect -2006 649218 -1974 649454
rect -1738 649218 -1654 649454
rect -1418 649218 -1386 649454
rect -2006 649134 -1386 649218
rect -2006 648898 -1974 649134
rect -1738 648898 -1654 649134
rect -1418 648898 -1386 649134
rect -2006 615454 -1386 648898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 581454 -1386 614898
rect -2006 581218 -1974 581454
rect -1738 581218 -1654 581454
rect -1418 581218 -1386 581454
rect -2006 581134 -1386 581218
rect -2006 580898 -1974 581134
rect -1738 580898 -1654 581134
rect -1418 580898 -1386 581134
rect -2006 547454 -1386 580898
rect -2006 547218 -1974 547454
rect -1738 547218 -1654 547454
rect -1418 547218 -1386 547454
rect -2006 547134 -1386 547218
rect -2006 546898 -1974 547134
rect -1738 546898 -1654 547134
rect -1418 546898 -1386 547134
rect -2006 513454 -1386 546898
rect -2006 513218 -1974 513454
rect -1738 513218 -1654 513454
rect -1418 513218 -1386 513454
rect -2006 513134 -1386 513218
rect -2006 512898 -1974 513134
rect -1738 512898 -1654 513134
rect -1418 512898 -1386 513134
rect -2006 479454 -1386 512898
rect -2006 479218 -1974 479454
rect -1738 479218 -1654 479454
rect -1418 479218 -1386 479454
rect -2006 479134 -1386 479218
rect -2006 478898 -1974 479134
rect -1738 478898 -1654 479134
rect -1418 478898 -1386 479134
rect -2006 445454 -1386 478898
rect -2006 445218 -1974 445454
rect -1738 445218 -1654 445454
rect -1418 445218 -1386 445454
rect -2006 445134 -1386 445218
rect -2006 444898 -1974 445134
rect -1738 444898 -1654 445134
rect -1418 444898 -1386 445134
rect -2006 411454 -1386 444898
rect -2006 411218 -1974 411454
rect -1738 411218 -1654 411454
rect -1418 411218 -1386 411454
rect -2006 411134 -1386 411218
rect -2006 410898 -1974 411134
rect -1738 410898 -1654 411134
rect -1418 410898 -1386 411134
rect -2006 377454 -1386 410898
rect -2006 377218 -1974 377454
rect -1738 377218 -1654 377454
rect -1418 377218 -1386 377454
rect -2006 377134 -1386 377218
rect -2006 376898 -1974 377134
rect -1738 376898 -1654 377134
rect -1418 376898 -1386 377134
rect -2006 343454 -1386 376898
rect -2006 343218 -1974 343454
rect -1738 343218 -1654 343454
rect -1418 343218 -1386 343454
rect -2006 343134 -1386 343218
rect -2006 342898 -1974 343134
rect -1738 342898 -1654 343134
rect -1418 342898 -1386 343134
rect -2006 309454 -1386 342898
rect -2006 309218 -1974 309454
rect -1738 309218 -1654 309454
rect -1418 309218 -1386 309454
rect -2006 309134 -1386 309218
rect -2006 308898 -1974 309134
rect -1738 308898 -1654 309134
rect -1418 308898 -1386 309134
rect -2006 275454 -1386 308898
rect -2006 275218 -1974 275454
rect -1738 275218 -1654 275454
rect -1418 275218 -1386 275454
rect -2006 275134 -1386 275218
rect -2006 274898 -1974 275134
rect -1738 274898 -1654 275134
rect -1418 274898 -1386 275134
rect -2006 241454 -1386 274898
rect -2006 241218 -1974 241454
rect -1738 241218 -1654 241454
rect -1418 241218 -1386 241454
rect -2006 241134 -1386 241218
rect -2006 240898 -1974 241134
rect -1738 240898 -1654 241134
rect -1418 240898 -1386 241134
rect -2006 207454 -1386 240898
rect -2006 207218 -1974 207454
rect -1738 207218 -1654 207454
rect -1418 207218 -1386 207454
rect -2006 207134 -1386 207218
rect -2006 206898 -1974 207134
rect -1738 206898 -1654 207134
rect -1418 206898 -1386 207134
rect -2006 173454 -1386 206898
rect -2006 173218 -1974 173454
rect -1738 173218 -1654 173454
rect -1418 173218 -1386 173454
rect -2006 173134 -1386 173218
rect -2006 172898 -1974 173134
rect -1738 172898 -1654 173134
rect -1418 172898 -1386 173134
rect -2006 139454 -1386 172898
rect -2006 139218 -1974 139454
rect -1738 139218 -1654 139454
rect -1418 139218 -1386 139454
rect -2006 139134 -1386 139218
rect -2006 138898 -1974 139134
rect -1738 138898 -1654 139134
rect -1418 138898 -1386 139134
rect -2006 105454 -1386 138898
rect -2006 105218 -1974 105454
rect -1738 105218 -1654 105454
rect -1418 105218 -1386 105454
rect -2006 105134 -1386 105218
rect -2006 104898 -1974 105134
rect -1738 104898 -1654 105134
rect -1418 104898 -1386 105134
rect -2006 71454 -1386 104898
rect -2006 71218 -1974 71454
rect -1738 71218 -1654 71454
rect -1418 71218 -1386 71454
rect -2006 71134 -1386 71218
rect -2006 70898 -1974 71134
rect -1738 70898 -1654 71134
rect -1418 70898 -1386 71134
rect -2006 37454 -1386 70898
rect -2006 37218 -1974 37454
rect -1738 37218 -1654 37454
rect -1418 37218 -1386 37454
rect -2006 37134 -1386 37218
rect -2006 36898 -1974 37134
rect -1738 36898 -1654 37134
rect -1418 36898 -1386 37134
rect -2006 3454 -1386 36898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 683454 2414 704282
rect 1794 683218 1826 683454
rect 2062 683218 2146 683454
rect 2382 683218 2414 683454
rect 1794 683134 2414 683218
rect 1794 682898 1826 683134
rect 2062 682898 2146 683134
rect 2382 682898 2414 683134
rect 1794 649454 2414 682898
rect 1794 649218 1826 649454
rect 2062 649218 2146 649454
rect 2382 649218 2414 649454
rect 1794 649134 2414 649218
rect 1794 648898 1826 649134
rect 2062 648898 2146 649134
rect 2382 648898 2414 649134
rect 1794 615454 2414 648898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 581454 2414 614898
rect 1794 581218 1826 581454
rect 2062 581218 2146 581454
rect 2382 581218 2414 581454
rect 1794 581134 2414 581218
rect 1794 580898 1826 581134
rect 2062 580898 2146 581134
rect 2382 580898 2414 581134
rect 1794 547454 2414 580898
rect 1794 547218 1826 547454
rect 2062 547218 2146 547454
rect 2382 547218 2414 547454
rect 1794 547134 2414 547218
rect 1794 546898 1826 547134
rect 2062 546898 2146 547134
rect 2382 546898 2414 547134
rect 1794 513454 2414 546898
rect 1794 513218 1826 513454
rect 2062 513218 2146 513454
rect 2382 513218 2414 513454
rect 1794 513134 2414 513218
rect 1794 512898 1826 513134
rect 2062 512898 2146 513134
rect 2382 512898 2414 513134
rect 1794 479454 2414 512898
rect 1794 479218 1826 479454
rect 2062 479218 2146 479454
rect 2382 479218 2414 479454
rect 1794 479134 2414 479218
rect 1794 478898 1826 479134
rect 2062 478898 2146 479134
rect 2382 478898 2414 479134
rect 1794 445454 2414 478898
rect 1794 445218 1826 445454
rect 2062 445218 2146 445454
rect 2382 445218 2414 445454
rect 1794 445134 2414 445218
rect 1794 444898 1826 445134
rect 2062 444898 2146 445134
rect 2382 444898 2414 445134
rect 1794 411454 2414 444898
rect 1794 411218 1826 411454
rect 2062 411218 2146 411454
rect 2382 411218 2414 411454
rect 1794 411134 2414 411218
rect 1794 410898 1826 411134
rect 2062 410898 2146 411134
rect 2382 410898 2414 411134
rect 1794 377454 2414 410898
rect 1794 377218 1826 377454
rect 2062 377218 2146 377454
rect 2382 377218 2414 377454
rect 1794 377134 2414 377218
rect 1794 376898 1826 377134
rect 2062 376898 2146 377134
rect 2382 376898 2414 377134
rect 1794 343454 2414 376898
rect 1794 343218 1826 343454
rect 2062 343218 2146 343454
rect 2382 343218 2414 343454
rect 1794 343134 2414 343218
rect 1794 342898 1826 343134
rect 2062 342898 2146 343134
rect 2382 342898 2414 343134
rect 1794 309454 2414 342898
rect 1794 309218 1826 309454
rect 2062 309218 2146 309454
rect 2382 309218 2414 309454
rect 1794 309134 2414 309218
rect 1794 308898 1826 309134
rect 2062 308898 2146 309134
rect 2382 308898 2414 309134
rect 1794 275454 2414 308898
rect 1794 275218 1826 275454
rect 2062 275218 2146 275454
rect 2382 275218 2414 275454
rect 1794 275134 2414 275218
rect 1794 274898 1826 275134
rect 2062 274898 2146 275134
rect 2382 274898 2414 275134
rect 1794 241454 2414 274898
rect 1794 241218 1826 241454
rect 2062 241218 2146 241454
rect 2382 241218 2414 241454
rect 1794 241134 2414 241218
rect 1794 240898 1826 241134
rect 2062 240898 2146 241134
rect 2382 240898 2414 241134
rect 1794 207454 2414 240898
rect 1794 207218 1826 207454
rect 2062 207218 2146 207454
rect 2382 207218 2414 207454
rect 1794 207134 2414 207218
rect 1794 206898 1826 207134
rect 2062 206898 2146 207134
rect 2382 206898 2414 207134
rect 1794 173454 2414 206898
rect 1794 173218 1826 173454
rect 2062 173218 2146 173454
rect 2382 173218 2414 173454
rect 1794 173134 2414 173218
rect 1794 172898 1826 173134
rect 2062 172898 2146 173134
rect 2382 172898 2414 173134
rect 1794 139454 2414 172898
rect 1794 139218 1826 139454
rect 2062 139218 2146 139454
rect 2382 139218 2414 139454
rect 1794 139134 2414 139218
rect 1794 138898 1826 139134
rect 2062 138898 2146 139134
rect 2382 138898 2414 139134
rect 1794 105454 2414 138898
rect 1794 105218 1826 105454
rect 2062 105218 2146 105454
rect 2382 105218 2414 105454
rect 1794 105134 2414 105218
rect 1794 104898 1826 105134
rect 2062 104898 2146 105134
rect 2382 104898 2414 105134
rect 1794 71454 2414 104898
rect 1794 71218 1826 71454
rect 2062 71218 2146 71454
rect 2382 71218 2414 71454
rect 1794 71134 2414 71218
rect 1794 70898 1826 71134
rect 2062 70898 2146 71134
rect 2382 70898 2414 71134
rect 1794 37454 2414 70898
rect 1794 37218 1826 37454
rect 2062 37218 2146 37454
rect 2382 37218 2414 37454
rect 1794 37134 2414 37218
rect 1794 36898 1826 37134
rect 2062 36898 2146 37134
rect 2382 36898 2414 37134
rect 1794 3454 2414 36898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 687174 6134 705242
rect 5514 686938 5546 687174
rect 5782 686938 5866 687174
rect 6102 686938 6134 687174
rect 5514 686854 6134 686938
rect 5514 686618 5546 686854
rect 5782 686618 5866 686854
rect 6102 686618 6134 686854
rect 5514 653174 6134 686618
rect 5514 652938 5546 653174
rect 5782 652938 5866 653174
rect 6102 652938 6134 653174
rect 5514 652854 6134 652938
rect 5514 652618 5546 652854
rect 5782 652618 5866 652854
rect 6102 652618 6134 652854
rect 5514 619174 6134 652618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 585174 6134 618618
rect 5514 584938 5546 585174
rect 5782 584938 5866 585174
rect 6102 584938 6134 585174
rect 5514 584854 6134 584938
rect 5514 584618 5546 584854
rect 5782 584618 5866 584854
rect 6102 584618 6134 584854
rect 5514 551174 6134 584618
rect 5514 550938 5546 551174
rect 5782 550938 5866 551174
rect 6102 550938 6134 551174
rect 5514 550854 6134 550938
rect 5514 550618 5546 550854
rect 5782 550618 5866 550854
rect 6102 550618 6134 550854
rect 5514 517174 6134 550618
rect 5514 516938 5546 517174
rect 5782 516938 5866 517174
rect 6102 516938 6134 517174
rect 5514 516854 6134 516938
rect 5514 516618 5546 516854
rect 5782 516618 5866 516854
rect 6102 516618 6134 516854
rect 5514 483174 6134 516618
rect 5514 482938 5546 483174
rect 5782 482938 5866 483174
rect 6102 482938 6134 483174
rect 5514 482854 6134 482938
rect 5514 482618 5546 482854
rect 5782 482618 5866 482854
rect 6102 482618 6134 482854
rect 5514 449174 6134 482618
rect 5514 448938 5546 449174
rect 5782 448938 5866 449174
rect 6102 448938 6134 449174
rect 5514 448854 6134 448938
rect 5514 448618 5546 448854
rect 5782 448618 5866 448854
rect 6102 448618 6134 448854
rect 5514 415174 6134 448618
rect 5514 414938 5546 415174
rect 5782 414938 5866 415174
rect 6102 414938 6134 415174
rect 5514 414854 6134 414938
rect 5514 414618 5546 414854
rect 5782 414618 5866 414854
rect 6102 414618 6134 414854
rect 5514 381174 6134 414618
rect 5514 380938 5546 381174
rect 5782 380938 5866 381174
rect 6102 380938 6134 381174
rect 5514 380854 6134 380938
rect 5514 380618 5546 380854
rect 5782 380618 5866 380854
rect 6102 380618 6134 380854
rect 5514 347174 6134 380618
rect 5514 346938 5546 347174
rect 5782 346938 5866 347174
rect 6102 346938 6134 347174
rect 5514 346854 6134 346938
rect 5514 346618 5546 346854
rect 5782 346618 5866 346854
rect 6102 346618 6134 346854
rect 5514 313174 6134 346618
rect 5514 312938 5546 313174
rect 5782 312938 5866 313174
rect 6102 312938 6134 313174
rect 5514 312854 6134 312938
rect 5514 312618 5546 312854
rect 5782 312618 5866 312854
rect 6102 312618 6134 312854
rect 5514 279174 6134 312618
rect 5514 278938 5546 279174
rect 5782 278938 5866 279174
rect 6102 278938 6134 279174
rect 5514 278854 6134 278938
rect 5514 278618 5546 278854
rect 5782 278618 5866 278854
rect 6102 278618 6134 278854
rect 5514 245174 6134 278618
rect 5514 244938 5546 245174
rect 5782 244938 5866 245174
rect 6102 244938 6134 245174
rect 5514 244854 6134 244938
rect 5514 244618 5546 244854
rect 5782 244618 5866 244854
rect 6102 244618 6134 244854
rect 5514 211174 6134 244618
rect 5514 210938 5546 211174
rect 5782 210938 5866 211174
rect 6102 210938 6134 211174
rect 5514 210854 6134 210938
rect 5514 210618 5546 210854
rect 5782 210618 5866 210854
rect 6102 210618 6134 210854
rect 5514 177174 6134 210618
rect 5514 176938 5546 177174
rect 5782 176938 5866 177174
rect 6102 176938 6134 177174
rect 5514 176854 6134 176938
rect 5514 176618 5546 176854
rect 5782 176618 5866 176854
rect 6102 176618 6134 176854
rect 5514 143174 6134 176618
rect 5514 142938 5546 143174
rect 5782 142938 5866 143174
rect 6102 142938 6134 143174
rect 5514 142854 6134 142938
rect 5514 142618 5546 142854
rect 5782 142618 5866 142854
rect 6102 142618 6134 142854
rect 5514 109174 6134 142618
rect 5514 108938 5546 109174
rect 5782 108938 5866 109174
rect 6102 108938 6134 109174
rect 5514 108854 6134 108938
rect 5514 108618 5546 108854
rect 5782 108618 5866 108854
rect 6102 108618 6134 108854
rect 5514 75174 6134 108618
rect 5514 74938 5546 75174
rect 5782 74938 5866 75174
rect 6102 74938 6134 75174
rect 5514 74854 6134 74938
rect 5514 74618 5546 74854
rect 5782 74618 5866 74854
rect 6102 74618 6134 74854
rect 5514 41174 6134 74618
rect 5514 40938 5546 41174
rect 5782 40938 5866 41174
rect 6102 40938 6134 41174
rect 5514 40854 6134 40938
rect 5514 40618 5546 40854
rect 5782 40618 5866 40854
rect 6102 40618 6134 40854
rect 5514 7174 6134 40618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 690894 9854 706202
rect 9234 690658 9266 690894
rect 9502 690658 9586 690894
rect 9822 690658 9854 690894
rect 9234 690574 9854 690658
rect 9234 690338 9266 690574
rect 9502 690338 9586 690574
rect 9822 690338 9854 690574
rect 9234 656894 9854 690338
rect 9234 656658 9266 656894
rect 9502 656658 9586 656894
rect 9822 656658 9854 656894
rect 9234 656574 9854 656658
rect 9234 656338 9266 656574
rect 9502 656338 9586 656574
rect 9822 656338 9854 656574
rect 9234 622894 9854 656338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 588894 9854 622338
rect 9234 588658 9266 588894
rect 9502 588658 9586 588894
rect 9822 588658 9854 588894
rect 9234 588574 9854 588658
rect 9234 588338 9266 588574
rect 9502 588338 9586 588574
rect 9822 588338 9854 588574
rect 9234 554894 9854 588338
rect 9234 554658 9266 554894
rect 9502 554658 9586 554894
rect 9822 554658 9854 554894
rect 9234 554574 9854 554658
rect 9234 554338 9266 554574
rect 9502 554338 9586 554574
rect 9822 554338 9854 554574
rect 9234 520894 9854 554338
rect 9234 520658 9266 520894
rect 9502 520658 9586 520894
rect 9822 520658 9854 520894
rect 9234 520574 9854 520658
rect 9234 520338 9266 520574
rect 9502 520338 9586 520574
rect 9822 520338 9854 520574
rect 9234 486894 9854 520338
rect 9234 486658 9266 486894
rect 9502 486658 9586 486894
rect 9822 486658 9854 486894
rect 9234 486574 9854 486658
rect 9234 486338 9266 486574
rect 9502 486338 9586 486574
rect 9822 486338 9854 486574
rect 9234 452894 9854 486338
rect 9234 452658 9266 452894
rect 9502 452658 9586 452894
rect 9822 452658 9854 452894
rect 9234 452574 9854 452658
rect 9234 452338 9266 452574
rect 9502 452338 9586 452574
rect 9822 452338 9854 452574
rect 9234 418894 9854 452338
rect 9234 418658 9266 418894
rect 9502 418658 9586 418894
rect 9822 418658 9854 418894
rect 9234 418574 9854 418658
rect 9234 418338 9266 418574
rect 9502 418338 9586 418574
rect 9822 418338 9854 418574
rect 9234 384894 9854 418338
rect 9234 384658 9266 384894
rect 9502 384658 9586 384894
rect 9822 384658 9854 384894
rect 9234 384574 9854 384658
rect 9234 384338 9266 384574
rect 9502 384338 9586 384574
rect 9822 384338 9854 384574
rect 9234 350894 9854 384338
rect 9234 350658 9266 350894
rect 9502 350658 9586 350894
rect 9822 350658 9854 350894
rect 9234 350574 9854 350658
rect 9234 350338 9266 350574
rect 9502 350338 9586 350574
rect 9822 350338 9854 350574
rect 9234 316894 9854 350338
rect 9234 316658 9266 316894
rect 9502 316658 9586 316894
rect 9822 316658 9854 316894
rect 9234 316574 9854 316658
rect 9234 316338 9266 316574
rect 9502 316338 9586 316574
rect 9822 316338 9854 316574
rect 9234 282894 9854 316338
rect 9234 282658 9266 282894
rect 9502 282658 9586 282894
rect 9822 282658 9854 282894
rect 9234 282574 9854 282658
rect 9234 282338 9266 282574
rect 9502 282338 9586 282574
rect 9822 282338 9854 282574
rect 9234 248894 9854 282338
rect 9234 248658 9266 248894
rect 9502 248658 9586 248894
rect 9822 248658 9854 248894
rect 9234 248574 9854 248658
rect 9234 248338 9266 248574
rect 9502 248338 9586 248574
rect 9822 248338 9854 248574
rect 9234 214894 9854 248338
rect 9234 214658 9266 214894
rect 9502 214658 9586 214894
rect 9822 214658 9854 214894
rect 9234 214574 9854 214658
rect 9234 214338 9266 214574
rect 9502 214338 9586 214574
rect 9822 214338 9854 214574
rect 9234 180894 9854 214338
rect 9234 180658 9266 180894
rect 9502 180658 9586 180894
rect 9822 180658 9854 180894
rect 9234 180574 9854 180658
rect 9234 180338 9266 180574
rect 9502 180338 9586 180574
rect 9822 180338 9854 180574
rect 9234 146894 9854 180338
rect 9234 146658 9266 146894
rect 9502 146658 9586 146894
rect 9822 146658 9854 146894
rect 9234 146574 9854 146658
rect 9234 146338 9266 146574
rect 9502 146338 9586 146574
rect 9822 146338 9854 146574
rect 9234 112894 9854 146338
rect 9234 112658 9266 112894
rect 9502 112658 9586 112894
rect 9822 112658 9854 112894
rect 9234 112574 9854 112658
rect 9234 112338 9266 112574
rect 9502 112338 9586 112574
rect 9822 112338 9854 112574
rect 9234 78894 9854 112338
rect 9234 78658 9266 78894
rect 9502 78658 9586 78894
rect 9822 78658 9854 78894
rect 9234 78574 9854 78658
rect 9234 78338 9266 78574
rect 9502 78338 9586 78574
rect 9822 78338 9854 78574
rect 9234 44894 9854 78338
rect 9234 44658 9266 44894
rect 9502 44658 9586 44894
rect 9822 44658 9854 44894
rect 9234 44574 9854 44658
rect 9234 44338 9266 44574
rect 9502 44338 9586 44574
rect 9822 44338 9854 44574
rect 9234 10894 9854 44338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 694614 13574 707162
rect 12954 694378 12986 694614
rect 13222 694378 13306 694614
rect 13542 694378 13574 694614
rect 12954 694294 13574 694378
rect 12954 694058 12986 694294
rect 13222 694058 13306 694294
rect 13542 694058 13574 694294
rect 12954 660614 13574 694058
rect 12954 660378 12986 660614
rect 13222 660378 13306 660614
rect 13542 660378 13574 660614
rect 12954 660294 13574 660378
rect 12954 660058 12986 660294
rect 13222 660058 13306 660294
rect 13542 660058 13574 660294
rect 12954 626614 13574 660058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 592614 13574 626058
rect 12954 592378 12986 592614
rect 13222 592378 13306 592614
rect 13542 592378 13574 592614
rect 12954 592294 13574 592378
rect 12954 592058 12986 592294
rect 13222 592058 13306 592294
rect 13542 592058 13574 592294
rect 12954 558614 13574 592058
rect 12954 558378 12986 558614
rect 13222 558378 13306 558614
rect 13542 558378 13574 558614
rect 12954 558294 13574 558378
rect 12954 558058 12986 558294
rect 13222 558058 13306 558294
rect 13542 558058 13574 558294
rect 12954 524614 13574 558058
rect 12954 524378 12986 524614
rect 13222 524378 13306 524614
rect 13542 524378 13574 524614
rect 12954 524294 13574 524378
rect 12954 524058 12986 524294
rect 13222 524058 13306 524294
rect 13542 524058 13574 524294
rect 12954 490614 13574 524058
rect 12954 490378 12986 490614
rect 13222 490378 13306 490614
rect 13542 490378 13574 490614
rect 12954 490294 13574 490378
rect 12954 490058 12986 490294
rect 13222 490058 13306 490294
rect 13542 490058 13574 490294
rect 12954 456614 13574 490058
rect 12954 456378 12986 456614
rect 13222 456378 13306 456614
rect 13542 456378 13574 456614
rect 12954 456294 13574 456378
rect 12954 456058 12986 456294
rect 13222 456058 13306 456294
rect 13542 456058 13574 456294
rect 12954 422614 13574 456058
rect 12954 422378 12986 422614
rect 13222 422378 13306 422614
rect 13542 422378 13574 422614
rect 12954 422294 13574 422378
rect 12954 422058 12986 422294
rect 13222 422058 13306 422294
rect 13542 422058 13574 422294
rect 12954 388614 13574 422058
rect 12954 388378 12986 388614
rect 13222 388378 13306 388614
rect 13542 388378 13574 388614
rect 12954 388294 13574 388378
rect 12954 388058 12986 388294
rect 13222 388058 13306 388294
rect 13542 388058 13574 388294
rect 12954 354614 13574 388058
rect 12954 354378 12986 354614
rect 13222 354378 13306 354614
rect 13542 354378 13574 354614
rect 12954 354294 13574 354378
rect 12954 354058 12986 354294
rect 13222 354058 13306 354294
rect 13542 354058 13574 354294
rect 12954 320614 13574 354058
rect 12954 320378 12986 320614
rect 13222 320378 13306 320614
rect 13542 320378 13574 320614
rect 12954 320294 13574 320378
rect 12954 320058 12986 320294
rect 13222 320058 13306 320294
rect 13542 320058 13574 320294
rect 12954 286614 13574 320058
rect 12954 286378 12986 286614
rect 13222 286378 13306 286614
rect 13542 286378 13574 286614
rect 12954 286294 13574 286378
rect 12954 286058 12986 286294
rect 13222 286058 13306 286294
rect 13542 286058 13574 286294
rect 12954 252614 13574 286058
rect 12954 252378 12986 252614
rect 13222 252378 13306 252614
rect 13542 252378 13574 252614
rect 12954 252294 13574 252378
rect 12954 252058 12986 252294
rect 13222 252058 13306 252294
rect 13542 252058 13574 252294
rect 12954 218614 13574 252058
rect 12954 218378 12986 218614
rect 13222 218378 13306 218614
rect 13542 218378 13574 218614
rect 12954 218294 13574 218378
rect 12954 218058 12986 218294
rect 13222 218058 13306 218294
rect 13542 218058 13574 218294
rect 12954 184614 13574 218058
rect 12954 184378 12986 184614
rect 13222 184378 13306 184614
rect 13542 184378 13574 184614
rect 12954 184294 13574 184378
rect 12954 184058 12986 184294
rect 13222 184058 13306 184294
rect 13542 184058 13574 184294
rect 12954 150614 13574 184058
rect 12954 150378 12986 150614
rect 13222 150378 13306 150614
rect 13542 150378 13574 150614
rect 12954 150294 13574 150378
rect 12954 150058 12986 150294
rect 13222 150058 13306 150294
rect 13542 150058 13574 150294
rect 12954 116614 13574 150058
rect 12954 116378 12986 116614
rect 13222 116378 13306 116614
rect 13542 116378 13574 116614
rect 12954 116294 13574 116378
rect 12954 116058 12986 116294
rect 13222 116058 13306 116294
rect 13542 116058 13574 116294
rect 12954 82614 13574 116058
rect 12954 82378 12986 82614
rect 13222 82378 13306 82614
rect 13542 82378 13574 82614
rect 12954 82294 13574 82378
rect 12954 82058 12986 82294
rect 13222 82058 13306 82294
rect 13542 82058 13574 82294
rect 12954 48614 13574 82058
rect 12954 48378 12986 48614
rect 13222 48378 13306 48614
rect 13542 48378 13574 48614
rect 12954 48294 13574 48378
rect 12954 48058 12986 48294
rect 13222 48058 13306 48294
rect 13542 48058 13574 48294
rect 12954 14614 13574 48058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 698334 17294 708122
rect 16674 698098 16706 698334
rect 16942 698098 17026 698334
rect 17262 698098 17294 698334
rect 16674 698014 17294 698098
rect 16674 697778 16706 698014
rect 16942 697778 17026 698014
rect 17262 697778 17294 698014
rect 16674 664334 17294 697778
rect 16674 664098 16706 664334
rect 16942 664098 17026 664334
rect 17262 664098 17294 664334
rect 16674 664014 17294 664098
rect 16674 663778 16706 664014
rect 16942 663778 17026 664014
rect 17262 663778 17294 664014
rect 16674 630334 17294 663778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 596334 17294 629778
rect 16674 596098 16706 596334
rect 16942 596098 17026 596334
rect 17262 596098 17294 596334
rect 16674 596014 17294 596098
rect 16674 595778 16706 596014
rect 16942 595778 17026 596014
rect 17262 595778 17294 596014
rect 16674 562334 17294 595778
rect 16674 562098 16706 562334
rect 16942 562098 17026 562334
rect 17262 562098 17294 562334
rect 16674 562014 17294 562098
rect 16674 561778 16706 562014
rect 16942 561778 17026 562014
rect 17262 561778 17294 562014
rect 16674 528334 17294 561778
rect 16674 528098 16706 528334
rect 16942 528098 17026 528334
rect 17262 528098 17294 528334
rect 16674 528014 17294 528098
rect 16674 527778 16706 528014
rect 16942 527778 17026 528014
rect 17262 527778 17294 528014
rect 16674 494334 17294 527778
rect 16674 494098 16706 494334
rect 16942 494098 17026 494334
rect 17262 494098 17294 494334
rect 16674 494014 17294 494098
rect 16674 493778 16706 494014
rect 16942 493778 17026 494014
rect 17262 493778 17294 494014
rect 16674 460334 17294 493778
rect 16674 460098 16706 460334
rect 16942 460098 17026 460334
rect 17262 460098 17294 460334
rect 16674 460014 17294 460098
rect 16674 459778 16706 460014
rect 16942 459778 17026 460014
rect 17262 459778 17294 460014
rect 16674 426334 17294 459778
rect 16674 426098 16706 426334
rect 16942 426098 17026 426334
rect 17262 426098 17294 426334
rect 16674 426014 17294 426098
rect 16674 425778 16706 426014
rect 16942 425778 17026 426014
rect 17262 425778 17294 426014
rect 16674 392334 17294 425778
rect 16674 392098 16706 392334
rect 16942 392098 17026 392334
rect 17262 392098 17294 392334
rect 16674 392014 17294 392098
rect 16674 391778 16706 392014
rect 16942 391778 17026 392014
rect 17262 391778 17294 392014
rect 16674 358334 17294 391778
rect 16674 358098 16706 358334
rect 16942 358098 17026 358334
rect 17262 358098 17294 358334
rect 16674 358014 17294 358098
rect 16674 357778 16706 358014
rect 16942 357778 17026 358014
rect 17262 357778 17294 358014
rect 16674 324334 17294 357778
rect 16674 324098 16706 324334
rect 16942 324098 17026 324334
rect 17262 324098 17294 324334
rect 16674 324014 17294 324098
rect 16674 323778 16706 324014
rect 16942 323778 17026 324014
rect 17262 323778 17294 324014
rect 16674 290334 17294 323778
rect 16674 290098 16706 290334
rect 16942 290098 17026 290334
rect 17262 290098 17294 290334
rect 16674 290014 17294 290098
rect 16674 289778 16706 290014
rect 16942 289778 17026 290014
rect 17262 289778 17294 290014
rect 16674 256334 17294 289778
rect 16674 256098 16706 256334
rect 16942 256098 17026 256334
rect 17262 256098 17294 256334
rect 16674 256014 17294 256098
rect 16674 255778 16706 256014
rect 16942 255778 17026 256014
rect 17262 255778 17294 256014
rect 16674 222334 17294 255778
rect 16674 222098 16706 222334
rect 16942 222098 17026 222334
rect 17262 222098 17294 222334
rect 16674 222014 17294 222098
rect 16674 221778 16706 222014
rect 16942 221778 17026 222014
rect 17262 221778 17294 222014
rect 16674 188334 17294 221778
rect 16674 188098 16706 188334
rect 16942 188098 17026 188334
rect 17262 188098 17294 188334
rect 16674 188014 17294 188098
rect 16674 187778 16706 188014
rect 16942 187778 17026 188014
rect 17262 187778 17294 188014
rect 16674 154334 17294 187778
rect 16674 154098 16706 154334
rect 16942 154098 17026 154334
rect 17262 154098 17294 154334
rect 16674 154014 17294 154098
rect 16674 153778 16706 154014
rect 16942 153778 17026 154014
rect 17262 153778 17294 154014
rect 16674 120334 17294 153778
rect 16674 120098 16706 120334
rect 16942 120098 17026 120334
rect 17262 120098 17294 120334
rect 16674 120014 17294 120098
rect 16674 119778 16706 120014
rect 16942 119778 17026 120014
rect 17262 119778 17294 120014
rect 16674 86334 17294 119778
rect 16674 86098 16706 86334
rect 16942 86098 17026 86334
rect 17262 86098 17294 86334
rect 16674 86014 17294 86098
rect 16674 85778 16706 86014
rect 16942 85778 17026 86014
rect 17262 85778 17294 86014
rect 16674 52334 17294 85778
rect 16674 52098 16706 52334
rect 16942 52098 17026 52334
rect 17262 52098 17294 52334
rect 16674 52014 17294 52098
rect 16674 51778 16706 52014
rect 16942 51778 17026 52014
rect 17262 51778 17294 52014
rect 16674 18334 17294 51778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 668054 21014 709082
rect 20394 667818 20426 668054
rect 20662 667818 20746 668054
rect 20982 667818 21014 668054
rect 20394 667734 21014 667818
rect 20394 667498 20426 667734
rect 20662 667498 20746 667734
rect 20982 667498 21014 667734
rect 20394 634054 21014 667498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 600054 21014 633498
rect 20394 599818 20426 600054
rect 20662 599818 20746 600054
rect 20982 599818 21014 600054
rect 20394 599734 21014 599818
rect 20394 599498 20426 599734
rect 20662 599498 20746 599734
rect 20982 599498 21014 599734
rect 20394 566054 21014 599498
rect 20394 565818 20426 566054
rect 20662 565818 20746 566054
rect 20982 565818 21014 566054
rect 20394 565734 21014 565818
rect 20394 565498 20426 565734
rect 20662 565498 20746 565734
rect 20982 565498 21014 565734
rect 20394 532054 21014 565498
rect 20394 531818 20426 532054
rect 20662 531818 20746 532054
rect 20982 531818 21014 532054
rect 20394 531734 21014 531818
rect 20394 531498 20426 531734
rect 20662 531498 20746 531734
rect 20982 531498 21014 531734
rect 20394 498054 21014 531498
rect 20394 497818 20426 498054
rect 20662 497818 20746 498054
rect 20982 497818 21014 498054
rect 20394 497734 21014 497818
rect 20394 497498 20426 497734
rect 20662 497498 20746 497734
rect 20982 497498 21014 497734
rect 20394 464054 21014 497498
rect 20394 463818 20426 464054
rect 20662 463818 20746 464054
rect 20982 463818 21014 464054
rect 20394 463734 21014 463818
rect 20394 463498 20426 463734
rect 20662 463498 20746 463734
rect 20982 463498 21014 463734
rect 20394 430054 21014 463498
rect 20394 429818 20426 430054
rect 20662 429818 20746 430054
rect 20982 429818 21014 430054
rect 20394 429734 21014 429818
rect 20394 429498 20426 429734
rect 20662 429498 20746 429734
rect 20982 429498 21014 429734
rect 20394 396054 21014 429498
rect 20394 395818 20426 396054
rect 20662 395818 20746 396054
rect 20982 395818 21014 396054
rect 20394 395734 21014 395818
rect 20394 395498 20426 395734
rect 20662 395498 20746 395734
rect 20982 395498 21014 395734
rect 20394 362054 21014 395498
rect 20394 361818 20426 362054
rect 20662 361818 20746 362054
rect 20982 361818 21014 362054
rect 20394 361734 21014 361818
rect 20394 361498 20426 361734
rect 20662 361498 20746 361734
rect 20982 361498 21014 361734
rect 20394 328054 21014 361498
rect 20394 327818 20426 328054
rect 20662 327818 20746 328054
rect 20982 327818 21014 328054
rect 20394 327734 21014 327818
rect 20394 327498 20426 327734
rect 20662 327498 20746 327734
rect 20982 327498 21014 327734
rect 20394 294054 21014 327498
rect 20394 293818 20426 294054
rect 20662 293818 20746 294054
rect 20982 293818 21014 294054
rect 20394 293734 21014 293818
rect 20394 293498 20426 293734
rect 20662 293498 20746 293734
rect 20982 293498 21014 293734
rect 20394 260054 21014 293498
rect 20394 259818 20426 260054
rect 20662 259818 20746 260054
rect 20982 259818 21014 260054
rect 20394 259734 21014 259818
rect 20394 259498 20426 259734
rect 20662 259498 20746 259734
rect 20982 259498 21014 259734
rect 20394 226054 21014 259498
rect 20394 225818 20426 226054
rect 20662 225818 20746 226054
rect 20982 225818 21014 226054
rect 20394 225734 21014 225818
rect 20394 225498 20426 225734
rect 20662 225498 20746 225734
rect 20982 225498 21014 225734
rect 20394 192054 21014 225498
rect 20394 191818 20426 192054
rect 20662 191818 20746 192054
rect 20982 191818 21014 192054
rect 20394 191734 21014 191818
rect 20394 191498 20426 191734
rect 20662 191498 20746 191734
rect 20982 191498 21014 191734
rect 20394 158054 21014 191498
rect 20394 157818 20426 158054
rect 20662 157818 20746 158054
rect 20982 157818 21014 158054
rect 20394 157734 21014 157818
rect 20394 157498 20426 157734
rect 20662 157498 20746 157734
rect 20982 157498 21014 157734
rect 20394 124054 21014 157498
rect 20394 123818 20426 124054
rect 20662 123818 20746 124054
rect 20982 123818 21014 124054
rect 20394 123734 21014 123818
rect 20394 123498 20426 123734
rect 20662 123498 20746 123734
rect 20982 123498 21014 123734
rect 20394 90054 21014 123498
rect 20394 89818 20426 90054
rect 20662 89818 20746 90054
rect 20982 89818 21014 90054
rect 20394 89734 21014 89818
rect 20394 89498 20426 89734
rect 20662 89498 20746 89734
rect 20982 89498 21014 89734
rect 20394 56054 21014 89498
rect 20394 55818 20426 56054
rect 20662 55818 20746 56054
rect 20982 55818 21014 56054
rect 20394 55734 21014 55818
rect 20394 55498 20426 55734
rect 20662 55498 20746 55734
rect 20982 55498 21014 55734
rect 20394 22054 21014 55498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 671774 24734 710042
rect 24114 671538 24146 671774
rect 24382 671538 24466 671774
rect 24702 671538 24734 671774
rect 24114 671454 24734 671538
rect 24114 671218 24146 671454
rect 24382 671218 24466 671454
rect 24702 671218 24734 671454
rect 24114 637774 24734 671218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 603774 24734 637218
rect 24114 603538 24146 603774
rect 24382 603538 24466 603774
rect 24702 603538 24734 603774
rect 24114 603454 24734 603538
rect 24114 603218 24146 603454
rect 24382 603218 24466 603454
rect 24702 603218 24734 603454
rect 24114 569774 24734 603218
rect 24114 569538 24146 569774
rect 24382 569538 24466 569774
rect 24702 569538 24734 569774
rect 24114 569454 24734 569538
rect 24114 569218 24146 569454
rect 24382 569218 24466 569454
rect 24702 569218 24734 569454
rect 24114 535774 24734 569218
rect 24114 535538 24146 535774
rect 24382 535538 24466 535774
rect 24702 535538 24734 535774
rect 24114 535454 24734 535538
rect 24114 535218 24146 535454
rect 24382 535218 24466 535454
rect 24702 535218 24734 535454
rect 24114 501774 24734 535218
rect 24114 501538 24146 501774
rect 24382 501538 24466 501774
rect 24702 501538 24734 501774
rect 24114 501454 24734 501538
rect 24114 501218 24146 501454
rect 24382 501218 24466 501454
rect 24702 501218 24734 501454
rect 24114 467774 24734 501218
rect 24114 467538 24146 467774
rect 24382 467538 24466 467774
rect 24702 467538 24734 467774
rect 24114 467454 24734 467538
rect 24114 467218 24146 467454
rect 24382 467218 24466 467454
rect 24702 467218 24734 467454
rect 24114 433774 24734 467218
rect 24114 433538 24146 433774
rect 24382 433538 24466 433774
rect 24702 433538 24734 433774
rect 24114 433454 24734 433538
rect 24114 433218 24146 433454
rect 24382 433218 24466 433454
rect 24702 433218 24734 433454
rect 24114 399774 24734 433218
rect 24114 399538 24146 399774
rect 24382 399538 24466 399774
rect 24702 399538 24734 399774
rect 24114 399454 24734 399538
rect 24114 399218 24146 399454
rect 24382 399218 24466 399454
rect 24702 399218 24734 399454
rect 24114 365774 24734 399218
rect 24114 365538 24146 365774
rect 24382 365538 24466 365774
rect 24702 365538 24734 365774
rect 24114 365454 24734 365538
rect 24114 365218 24146 365454
rect 24382 365218 24466 365454
rect 24702 365218 24734 365454
rect 24114 331774 24734 365218
rect 24114 331538 24146 331774
rect 24382 331538 24466 331774
rect 24702 331538 24734 331774
rect 24114 331454 24734 331538
rect 24114 331218 24146 331454
rect 24382 331218 24466 331454
rect 24702 331218 24734 331454
rect 24114 297774 24734 331218
rect 24114 297538 24146 297774
rect 24382 297538 24466 297774
rect 24702 297538 24734 297774
rect 24114 297454 24734 297538
rect 24114 297218 24146 297454
rect 24382 297218 24466 297454
rect 24702 297218 24734 297454
rect 24114 263774 24734 297218
rect 24114 263538 24146 263774
rect 24382 263538 24466 263774
rect 24702 263538 24734 263774
rect 24114 263454 24734 263538
rect 24114 263218 24146 263454
rect 24382 263218 24466 263454
rect 24702 263218 24734 263454
rect 24114 229774 24734 263218
rect 24114 229538 24146 229774
rect 24382 229538 24466 229774
rect 24702 229538 24734 229774
rect 24114 229454 24734 229538
rect 24114 229218 24146 229454
rect 24382 229218 24466 229454
rect 24702 229218 24734 229454
rect 24114 195774 24734 229218
rect 24114 195538 24146 195774
rect 24382 195538 24466 195774
rect 24702 195538 24734 195774
rect 24114 195454 24734 195538
rect 24114 195218 24146 195454
rect 24382 195218 24466 195454
rect 24702 195218 24734 195454
rect 24114 161774 24734 195218
rect 24114 161538 24146 161774
rect 24382 161538 24466 161774
rect 24702 161538 24734 161774
rect 24114 161454 24734 161538
rect 24114 161218 24146 161454
rect 24382 161218 24466 161454
rect 24702 161218 24734 161454
rect 24114 127774 24734 161218
rect 24114 127538 24146 127774
rect 24382 127538 24466 127774
rect 24702 127538 24734 127774
rect 24114 127454 24734 127538
rect 24114 127218 24146 127454
rect 24382 127218 24466 127454
rect 24702 127218 24734 127454
rect 24114 93774 24734 127218
rect 24114 93538 24146 93774
rect 24382 93538 24466 93774
rect 24702 93538 24734 93774
rect 24114 93454 24734 93538
rect 24114 93218 24146 93454
rect 24382 93218 24466 93454
rect 24702 93218 24734 93454
rect 24114 59774 24734 93218
rect 24114 59538 24146 59774
rect 24382 59538 24466 59774
rect 24702 59538 24734 59774
rect 24114 59454 24734 59538
rect 24114 59218 24146 59454
rect 24382 59218 24466 59454
rect 24702 59218 24734 59454
rect 24114 25774 24734 59218
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 675494 28454 711002
rect 27834 675258 27866 675494
rect 28102 675258 28186 675494
rect 28422 675258 28454 675494
rect 27834 675174 28454 675258
rect 27834 674938 27866 675174
rect 28102 674938 28186 675174
rect 28422 674938 28454 675174
rect 27834 641494 28454 674938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 607494 28454 640938
rect 27834 607258 27866 607494
rect 28102 607258 28186 607494
rect 28422 607258 28454 607494
rect 27834 607174 28454 607258
rect 27834 606938 27866 607174
rect 28102 606938 28186 607174
rect 28422 606938 28454 607174
rect 27834 573494 28454 606938
rect 27834 573258 27866 573494
rect 28102 573258 28186 573494
rect 28422 573258 28454 573494
rect 27834 573174 28454 573258
rect 27834 572938 27866 573174
rect 28102 572938 28186 573174
rect 28422 572938 28454 573174
rect 27834 539494 28454 572938
rect 27834 539258 27866 539494
rect 28102 539258 28186 539494
rect 28422 539258 28454 539494
rect 27834 539174 28454 539258
rect 27834 538938 27866 539174
rect 28102 538938 28186 539174
rect 28422 538938 28454 539174
rect 27834 505494 28454 538938
rect 27834 505258 27866 505494
rect 28102 505258 28186 505494
rect 28422 505258 28454 505494
rect 27834 505174 28454 505258
rect 27834 504938 27866 505174
rect 28102 504938 28186 505174
rect 28422 504938 28454 505174
rect 27834 471494 28454 504938
rect 27834 471258 27866 471494
rect 28102 471258 28186 471494
rect 28422 471258 28454 471494
rect 27834 471174 28454 471258
rect 27834 470938 27866 471174
rect 28102 470938 28186 471174
rect 28422 470938 28454 471174
rect 27834 437494 28454 470938
rect 27834 437258 27866 437494
rect 28102 437258 28186 437494
rect 28422 437258 28454 437494
rect 27834 437174 28454 437258
rect 27834 436938 27866 437174
rect 28102 436938 28186 437174
rect 28422 436938 28454 437174
rect 27834 403494 28454 436938
rect 27834 403258 27866 403494
rect 28102 403258 28186 403494
rect 28422 403258 28454 403494
rect 27834 403174 28454 403258
rect 27834 402938 27866 403174
rect 28102 402938 28186 403174
rect 28422 402938 28454 403174
rect 27834 369494 28454 402938
rect 27834 369258 27866 369494
rect 28102 369258 28186 369494
rect 28422 369258 28454 369494
rect 27834 369174 28454 369258
rect 27834 368938 27866 369174
rect 28102 368938 28186 369174
rect 28422 368938 28454 369174
rect 27834 335494 28454 368938
rect 27834 335258 27866 335494
rect 28102 335258 28186 335494
rect 28422 335258 28454 335494
rect 27834 335174 28454 335258
rect 27834 334938 27866 335174
rect 28102 334938 28186 335174
rect 28422 334938 28454 335174
rect 27834 301494 28454 334938
rect 27834 301258 27866 301494
rect 28102 301258 28186 301494
rect 28422 301258 28454 301494
rect 27834 301174 28454 301258
rect 27834 300938 27866 301174
rect 28102 300938 28186 301174
rect 28422 300938 28454 301174
rect 27834 267494 28454 300938
rect 27834 267258 27866 267494
rect 28102 267258 28186 267494
rect 28422 267258 28454 267494
rect 27834 267174 28454 267258
rect 27834 266938 27866 267174
rect 28102 266938 28186 267174
rect 28422 266938 28454 267174
rect 27834 233494 28454 266938
rect 27834 233258 27866 233494
rect 28102 233258 28186 233494
rect 28422 233258 28454 233494
rect 27834 233174 28454 233258
rect 27834 232938 27866 233174
rect 28102 232938 28186 233174
rect 28422 232938 28454 233174
rect 27834 199494 28454 232938
rect 27834 199258 27866 199494
rect 28102 199258 28186 199494
rect 28422 199258 28454 199494
rect 27834 199174 28454 199258
rect 27834 198938 27866 199174
rect 28102 198938 28186 199174
rect 28422 198938 28454 199174
rect 27834 165494 28454 198938
rect 27834 165258 27866 165494
rect 28102 165258 28186 165494
rect 28422 165258 28454 165494
rect 27834 165174 28454 165258
rect 27834 164938 27866 165174
rect 28102 164938 28186 165174
rect 28422 164938 28454 165174
rect 27834 131494 28454 164938
rect 27834 131258 27866 131494
rect 28102 131258 28186 131494
rect 28422 131258 28454 131494
rect 27834 131174 28454 131258
rect 27834 130938 27866 131174
rect 28102 130938 28186 131174
rect 28422 130938 28454 131174
rect 27834 97494 28454 130938
rect 27834 97258 27866 97494
rect 28102 97258 28186 97494
rect 28422 97258 28454 97494
rect 27834 97174 28454 97258
rect 27834 96938 27866 97174
rect 28102 96938 28186 97174
rect 28422 96938 28454 97174
rect 27834 63494 28454 96938
rect 27834 63258 27866 63494
rect 28102 63258 28186 63494
rect 28422 63258 28454 63494
rect 27834 63174 28454 63258
rect 27834 62938 27866 63174
rect 28102 62938 28186 63174
rect 28422 62938 28454 63174
rect 27834 29494 28454 62938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 35794 704838 36414 711590
rect 35794 704602 35826 704838
rect 36062 704602 36146 704838
rect 36382 704602 36414 704838
rect 35794 704518 36414 704602
rect 35794 704282 35826 704518
rect 36062 704282 36146 704518
rect 36382 704282 36414 704518
rect 35794 683454 36414 704282
rect 35794 683218 35826 683454
rect 36062 683218 36146 683454
rect 36382 683218 36414 683454
rect 35794 683134 36414 683218
rect 35794 682898 35826 683134
rect 36062 682898 36146 683134
rect 36382 682898 36414 683134
rect 35794 649454 36414 682898
rect 35794 649218 35826 649454
rect 36062 649218 36146 649454
rect 36382 649218 36414 649454
rect 35794 649134 36414 649218
rect 35794 648898 35826 649134
rect 36062 648898 36146 649134
rect 36382 648898 36414 649134
rect 35794 615454 36414 648898
rect 35794 615218 35826 615454
rect 36062 615218 36146 615454
rect 36382 615218 36414 615454
rect 35794 615134 36414 615218
rect 35794 614898 35826 615134
rect 36062 614898 36146 615134
rect 36382 614898 36414 615134
rect 35794 581454 36414 614898
rect 35794 581218 35826 581454
rect 36062 581218 36146 581454
rect 36382 581218 36414 581454
rect 35794 581134 36414 581218
rect 35794 580898 35826 581134
rect 36062 580898 36146 581134
rect 36382 580898 36414 581134
rect 35794 547454 36414 580898
rect 35794 547218 35826 547454
rect 36062 547218 36146 547454
rect 36382 547218 36414 547454
rect 35794 547134 36414 547218
rect 35794 546898 35826 547134
rect 36062 546898 36146 547134
rect 36382 546898 36414 547134
rect 35794 513454 36414 546898
rect 35794 513218 35826 513454
rect 36062 513218 36146 513454
rect 36382 513218 36414 513454
rect 35794 513134 36414 513218
rect 35794 512898 35826 513134
rect 36062 512898 36146 513134
rect 36382 512898 36414 513134
rect 35794 479454 36414 512898
rect 35794 479218 35826 479454
rect 36062 479218 36146 479454
rect 36382 479218 36414 479454
rect 35794 479134 36414 479218
rect 35794 478898 35826 479134
rect 36062 478898 36146 479134
rect 36382 478898 36414 479134
rect 35794 445454 36414 478898
rect 35794 445218 35826 445454
rect 36062 445218 36146 445454
rect 36382 445218 36414 445454
rect 35794 445134 36414 445218
rect 35794 444898 35826 445134
rect 36062 444898 36146 445134
rect 36382 444898 36414 445134
rect 35794 411454 36414 444898
rect 35794 411218 35826 411454
rect 36062 411218 36146 411454
rect 36382 411218 36414 411454
rect 35794 411134 36414 411218
rect 35794 410898 35826 411134
rect 36062 410898 36146 411134
rect 36382 410898 36414 411134
rect 35794 377454 36414 410898
rect 35794 377218 35826 377454
rect 36062 377218 36146 377454
rect 36382 377218 36414 377454
rect 35794 377134 36414 377218
rect 35794 376898 35826 377134
rect 36062 376898 36146 377134
rect 36382 376898 36414 377134
rect 35794 343454 36414 376898
rect 35794 343218 35826 343454
rect 36062 343218 36146 343454
rect 36382 343218 36414 343454
rect 35794 343134 36414 343218
rect 35794 342898 35826 343134
rect 36062 342898 36146 343134
rect 36382 342898 36414 343134
rect 35794 309454 36414 342898
rect 35794 309218 35826 309454
rect 36062 309218 36146 309454
rect 36382 309218 36414 309454
rect 35794 309134 36414 309218
rect 35794 308898 35826 309134
rect 36062 308898 36146 309134
rect 36382 308898 36414 309134
rect 35794 275454 36414 308898
rect 35794 275218 35826 275454
rect 36062 275218 36146 275454
rect 36382 275218 36414 275454
rect 35794 275134 36414 275218
rect 35794 274898 35826 275134
rect 36062 274898 36146 275134
rect 36382 274898 36414 275134
rect 35794 241454 36414 274898
rect 35794 241218 35826 241454
rect 36062 241218 36146 241454
rect 36382 241218 36414 241454
rect 35794 241134 36414 241218
rect 35794 240898 35826 241134
rect 36062 240898 36146 241134
rect 36382 240898 36414 241134
rect 35794 207454 36414 240898
rect 35794 207218 35826 207454
rect 36062 207218 36146 207454
rect 36382 207218 36414 207454
rect 35794 207134 36414 207218
rect 35794 206898 35826 207134
rect 36062 206898 36146 207134
rect 36382 206898 36414 207134
rect 35794 173454 36414 206898
rect 35794 173218 35826 173454
rect 36062 173218 36146 173454
rect 36382 173218 36414 173454
rect 35794 173134 36414 173218
rect 35794 172898 35826 173134
rect 36062 172898 36146 173134
rect 36382 172898 36414 173134
rect 35794 139454 36414 172898
rect 35794 139218 35826 139454
rect 36062 139218 36146 139454
rect 36382 139218 36414 139454
rect 35794 139134 36414 139218
rect 35794 138898 35826 139134
rect 36062 138898 36146 139134
rect 36382 138898 36414 139134
rect 35794 105454 36414 138898
rect 35794 105218 35826 105454
rect 36062 105218 36146 105454
rect 36382 105218 36414 105454
rect 35794 105134 36414 105218
rect 35794 104898 35826 105134
rect 36062 104898 36146 105134
rect 36382 104898 36414 105134
rect 35794 71454 36414 104898
rect 35794 71218 35826 71454
rect 36062 71218 36146 71454
rect 36382 71218 36414 71454
rect 35794 71134 36414 71218
rect 35794 70898 35826 71134
rect 36062 70898 36146 71134
rect 36382 70898 36414 71134
rect 35794 37454 36414 70898
rect 35794 37218 35826 37454
rect 36062 37218 36146 37454
rect 36382 37218 36414 37454
rect 35794 37134 36414 37218
rect 35794 36898 35826 37134
rect 36062 36898 36146 37134
rect 36382 36898 36414 37134
rect 35794 3454 36414 36898
rect 35794 3218 35826 3454
rect 36062 3218 36146 3454
rect 36382 3218 36414 3454
rect 35794 3134 36414 3218
rect 35794 2898 35826 3134
rect 36062 2898 36146 3134
rect 36382 2898 36414 3134
rect 35794 -346 36414 2898
rect 35794 -582 35826 -346
rect 36062 -582 36146 -346
rect 36382 -582 36414 -346
rect 35794 -666 36414 -582
rect 35794 -902 35826 -666
rect 36062 -902 36146 -666
rect 36382 -902 36414 -666
rect 35794 -7654 36414 -902
rect 39514 705798 40134 711590
rect 39514 705562 39546 705798
rect 39782 705562 39866 705798
rect 40102 705562 40134 705798
rect 39514 705478 40134 705562
rect 39514 705242 39546 705478
rect 39782 705242 39866 705478
rect 40102 705242 40134 705478
rect 39514 687174 40134 705242
rect 39514 686938 39546 687174
rect 39782 686938 39866 687174
rect 40102 686938 40134 687174
rect 39514 686854 40134 686938
rect 39514 686618 39546 686854
rect 39782 686618 39866 686854
rect 40102 686618 40134 686854
rect 39514 653174 40134 686618
rect 39514 652938 39546 653174
rect 39782 652938 39866 653174
rect 40102 652938 40134 653174
rect 39514 652854 40134 652938
rect 39514 652618 39546 652854
rect 39782 652618 39866 652854
rect 40102 652618 40134 652854
rect 39514 619174 40134 652618
rect 39514 618938 39546 619174
rect 39782 618938 39866 619174
rect 40102 618938 40134 619174
rect 39514 618854 40134 618938
rect 39514 618618 39546 618854
rect 39782 618618 39866 618854
rect 40102 618618 40134 618854
rect 39514 585174 40134 618618
rect 39514 584938 39546 585174
rect 39782 584938 39866 585174
rect 40102 584938 40134 585174
rect 39514 584854 40134 584938
rect 39514 584618 39546 584854
rect 39782 584618 39866 584854
rect 40102 584618 40134 584854
rect 39514 551174 40134 584618
rect 39514 550938 39546 551174
rect 39782 550938 39866 551174
rect 40102 550938 40134 551174
rect 39514 550854 40134 550938
rect 39514 550618 39546 550854
rect 39782 550618 39866 550854
rect 40102 550618 40134 550854
rect 39514 517174 40134 550618
rect 39514 516938 39546 517174
rect 39782 516938 39866 517174
rect 40102 516938 40134 517174
rect 39514 516854 40134 516938
rect 39514 516618 39546 516854
rect 39782 516618 39866 516854
rect 40102 516618 40134 516854
rect 39514 483174 40134 516618
rect 39514 482938 39546 483174
rect 39782 482938 39866 483174
rect 40102 482938 40134 483174
rect 39514 482854 40134 482938
rect 39514 482618 39546 482854
rect 39782 482618 39866 482854
rect 40102 482618 40134 482854
rect 39514 449174 40134 482618
rect 39514 448938 39546 449174
rect 39782 448938 39866 449174
rect 40102 448938 40134 449174
rect 39514 448854 40134 448938
rect 39514 448618 39546 448854
rect 39782 448618 39866 448854
rect 40102 448618 40134 448854
rect 39514 415174 40134 448618
rect 39514 414938 39546 415174
rect 39782 414938 39866 415174
rect 40102 414938 40134 415174
rect 39514 414854 40134 414938
rect 39514 414618 39546 414854
rect 39782 414618 39866 414854
rect 40102 414618 40134 414854
rect 39514 381174 40134 414618
rect 39514 380938 39546 381174
rect 39782 380938 39866 381174
rect 40102 380938 40134 381174
rect 39514 380854 40134 380938
rect 39514 380618 39546 380854
rect 39782 380618 39866 380854
rect 40102 380618 40134 380854
rect 39514 347174 40134 380618
rect 39514 346938 39546 347174
rect 39782 346938 39866 347174
rect 40102 346938 40134 347174
rect 39514 346854 40134 346938
rect 39514 346618 39546 346854
rect 39782 346618 39866 346854
rect 40102 346618 40134 346854
rect 39514 313174 40134 346618
rect 39514 312938 39546 313174
rect 39782 312938 39866 313174
rect 40102 312938 40134 313174
rect 39514 312854 40134 312938
rect 39514 312618 39546 312854
rect 39782 312618 39866 312854
rect 40102 312618 40134 312854
rect 39514 279174 40134 312618
rect 39514 278938 39546 279174
rect 39782 278938 39866 279174
rect 40102 278938 40134 279174
rect 39514 278854 40134 278938
rect 39514 278618 39546 278854
rect 39782 278618 39866 278854
rect 40102 278618 40134 278854
rect 39514 245174 40134 278618
rect 39514 244938 39546 245174
rect 39782 244938 39866 245174
rect 40102 244938 40134 245174
rect 39514 244854 40134 244938
rect 39514 244618 39546 244854
rect 39782 244618 39866 244854
rect 40102 244618 40134 244854
rect 39514 211174 40134 244618
rect 39514 210938 39546 211174
rect 39782 210938 39866 211174
rect 40102 210938 40134 211174
rect 39514 210854 40134 210938
rect 39514 210618 39546 210854
rect 39782 210618 39866 210854
rect 40102 210618 40134 210854
rect 39514 177174 40134 210618
rect 39514 176938 39546 177174
rect 39782 176938 39866 177174
rect 40102 176938 40134 177174
rect 39514 176854 40134 176938
rect 39514 176618 39546 176854
rect 39782 176618 39866 176854
rect 40102 176618 40134 176854
rect 39514 143174 40134 176618
rect 39514 142938 39546 143174
rect 39782 142938 39866 143174
rect 40102 142938 40134 143174
rect 39514 142854 40134 142938
rect 39514 142618 39546 142854
rect 39782 142618 39866 142854
rect 40102 142618 40134 142854
rect 39514 109174 40134 142618
rect 39514 108938 39546 109174
rect 39782 108938 39866 109174
rect 40102 108938 40134 109174
rect 39514 108854 40134 108938
rect 39514 108618 39546 108854
rect 39782 108618 39866 108854
rect 40102 108618 40134 108854
rect 39514 75174 40134 108618
rect 39514 74938 39546 75174
rect 39782 74938 39866 75174
rect 40102 74938 40134 75174
rect 39514 74854 40134 74938
rect 39514 74618 39546 74854
rect 39782 74618 39866 74854
rect 40102 74618 40134 74854
rect 39514 41174 40134 74618
rect 39514 40938 39546 41174
rect 39782 40938 39866 41174
rect 40102 40938 40134 41174
rect 39514 40854 40134 40938
rect 39514 40618 39546 40854
rect 39782 40618 39866 40854
rect 40102 40618 40134 40854
rect 39514 7174 40134 40618
rect 39514 6938 39546 7174
rect 39782 6938 39866 7174
rect 40102 6938 40134 7174
rect 39514 6854 40134 6938
rect 39514 6618 39546 6854
rect 39782 6618 39866 6854
rect 40102 6618 40134 6854
rect 39514 -1306 40134 6618
rect 39514 -1542 39546 -1306
rect 39782 -1542 39866 -1306
rect 40102 -1542 40134 -1306
rect 39514 -1626 40134 -1542
rect 39514 -1862 39546 -1626
rect 39782 -1862 39866 -1626
rect 40102 -1862 40134 -1626
rect 39514 -7654 40134 -1862
rect 43234 706758 43854 711590
rect 43234 706522 43266 706758
rect 43502 706522 43586 706758
rect 43822 706522 43854 706758
rect 43234 706438 43854 706522
rect 43234 706202 43266 706438
rect 43502 706202 43586 706438
rect 43822 706202 43854 706438
rect 43234 690894 43854 706202
rect 43234 690658 43266 690894
rect 43502 690658 43586 690894
rect 43822 690658 43854 690894
rect 43234 690574 43854 690658
rect 43234 690338 43266 690574
rect 43502 690338 43586 690574
rect 43822 690338 43854 690574
rect 43234 656894 43854 690338
rect 43234 656658 43266 656894
rect 43502 656658 43586 656894
rect 43822 656658 43854 656894
rect 43234 656574 43854 656658
rect 43234 656338 43266 656574
rect 43502 656338 43586 656574
rect 43822 656338 43854 656574
rect 43234 622894 43854 656338
rect 43234 622658 43266 622894
rect 43502 622658 43586 622894
rect 43822 622658 43854 622894
rect 43234 622574 43854 622658
rect 43234 622338 43266 622574
rect 43502 622338 43586 622574
rect 43822 622338 43854 622574
rect 43234 588894 43854 622338
rect 43234 588658 43266 588894
rect 43502 588658 43586 588894
rect 43822 588658 43854 588894
rect 43234 588574 43854 588658
rect 43234 588338 43266 588574
rect 43502 588338 43586 588574
rect 43822 588338 43854 588574
rect 43234 554894 43854 588338
rect 43234 554658 43266 554894
rect 43502 554658 43586 554894
rect 43822 554658 43854 554894
rect 43234 554574 43854 554658
rect 43234 554338 43266 554574
rect 43502 554338 43586 554574
rect 43822 554338 43854 554574
rect 43234 520894 43854 554338
rect 43234 520658 43266 520894
rect 43502 520658 43586 520894
rect 43822 520658 43854 520894
rect 43234 520574 43854 520658
rect 43234 520338 43266 520574
rect 43502 520338 43586 520574
rect 43822 520338 43854 520574
rect 43234 486894 43854 520338
rect 43234 486658 43266 486894
rect 43502 486658 43586 486894
rect 43822 486658 43854 486894
rect 43234 486574 43854 486658
rect 43234 486338 43266 486574
rect 43502 486338 43586 486574
rect 43822 486338 43854 486574
rect 43234 452894 43854 486338
rect 43234 452658 43266 452894
rect 43502 452658 43586 452894
rect 43822 452658 43854 452894
rect 43234 452574 43854 452658
rect 43234 452338 43266 452574
rect 43502 452338 43586 452574
rect 43822 452338 43854 452574
rect 43234 418894 43854 452338
rect 43234 418658 43266 418894
rect 43502 418658 43586 418894
rect 43822 418658 43854 418894
rect 43234 418574 43854 418658
rect 43234 418338 43266 418574
rect 43502 418338 43586 418574
rect 43822 418338 43854 418574
rect 43234 384894 43854 418338
rect 43234 384658 43266 384894
rect 43502 384658 43586 384894
rect 43822 384658 43854 384894
rect 43234 384574 43854 384658
rect 43234 384338 43266 384574
rect 43502 384338 43586 384574
rect 43822 384338 43854 384574
rect 43234 350894 43854 384338
rect 43234 350658 43266 350894
rect 43502 350658 43586 350894
rect 43822 350658 43854 350894
rect 43234 350574 43854 350658
rect 43234 350338 43266 350574
rect 43502 350338 43586 350574
rect 43822 350338 43854 350574
rect 43234 316894 43854 350338
rect 43234 316658 43266 316894
rect 43502 316658 43586 316894
rect 43822 316658 43854 316894
rect 43234 316574 43854 316658
rect 43234 316338 43266 316574
rect 43502 316338 43586 316574
rect 43822 316338 43854 316574
rect 43234 282894 43854 316338
rect 43234 282658 43266 282894
rect 43502 282658 43586 282894
rect 43822 282658 43854 282894
rect 43234 282574 43854 282658
rect 43234 282338 43266 282574
rect 43502 282338 43586 282574
rect 43822 282338 43854 282574
rect 43234 248894 43854 282338
rect 43234 248658 43266 248894
rect 43502 248658 43586 248894
rect 43822 248658 43854 248894
rect 43234 248574 43854 248658
rect 43234 248338 43266 248574
rect 43502 248338 43586 248574
rect 43822 248338 43854 248574
rect 43234 214894 43854 248338
rect 46954 707718 47574 711590
rect 46954 707482 46986 707718
rect 47222 707482 47306 707718
rect 47542 707482 47574 707718
rect 46954 707398 47574 707482
rect 46954 707162 46986 707398
rect 47222 707162 47306 707398
rect 47542 707162 47574 707398
rect 46954 694614 47574 707162
rect 46954 694378 46986 694614
rect 47222 694378 47306 694614
rect 47542 694378 47574 694614
rect 46954 694294 47574 694378
rect 46954 694058 46986 694294
rect 47222 694058 47306 694294
rect 47542 694058 47574 694294
rect 46954 660614 47574 694058
rect 46954 660378 46986 660614
rect 47222 660378 47306 660614
rect 47542 660378 47574 660614
rect 46954 660294 47574 660378
rect 46954 660058 46986 660294
rect 47222 660058 47306 660294
rect 47542 660058 47574 660294
rect 46954 626614 47574 660058
rect 46954 626378 46986 626614
rect 47222 626378 47306 626614
rect 47542 626378 47574 626614
rect 46954 626294 47574 626378
rect 46954 626058 46986 626294
rect 47222 626058 47306 626294
rect 47542 626058 47574 626294
rect 46954 592614 47574 626058
rect 46954 592378 46986 592614
rect 47222 592378 47306 592614
rect 47542 592378 47574 592614
rect 46954 592294 47574 592378
rect 46954 592058 46986 592294
rect 47222 592058 47306 592294
rect 47542 592058 47574 592294
rect 46954 558614 47574 592058
rect 46954 558378 46986 558614
rect 47222 558378 47306 558614
rect 47542 558378 47574 558614
rect 46954 558294 47574 558378
rect 46954 558058 46986 558294
rect 47222 558058 47306 558294
rect 47542 558058 47574 558294
rect 46954 524614 47574 558058
rect 46954 524378 46986 524614
rect 47222 524378 47306 524614
rect 47542 524378 47574 524614
rect 46954 524294 47574 524378
rect 46954 524058 46986 524294
rect 47222 524058 47306 524294
rect 47542 524058 47574 524294
rect 46954 490614 47574 524058
rect 46954 490378 46986 490614
rect 47222 490378 47306 490614
rect 47542 490378 47574 490614
rect 46954 490294 47574 490378
rect 46954 490058 46986 490294
rect 47222 490058 47306 490294
rect 47542 490058 47574 490294
rect 46954 456614 47574 490058
rect 46954 456378 46986 456614
rect 47222 456378 47306 456614
rect 47542 456378 47574 456614
rect 46954 456294 47574 456378
rect 46954 456058 46986 456294
rect 47222 456058 47306 456294
rect 47542 456058 47574 456294
rect 46954 422614 47574 456058
rect 46954 422378 46986 422614
rect 47222 422378 47306 422614
rect 47542 422378 47574 422614
rect 46954 422294 47574 422378
rect 46954 422058 46986 422294
rect 47222 422058 47306 422294
rect 47542 422058 47574 422294
rect 46954 388614 47574 422058
rect 46954 388378 46986 388614
rect 47222 388378 47306 388614
rect 47542 388378 47574 388614
rect 46954 388294 47574 388378
rect 46954 388058 46986 388294
rect 47222 388058 47306 388294
rect 47542 388058 47574 388294
rect 46954 354614 47574 388058
rect 46954 354378 46986 354614
rect 47222 354378 47306 354614
rect 47542 354378 47574 354614
rect 46954 354294 47574 354378
rect 46954 354058 46986 354294
rect 47222 354058 47306 354294
rect 47542 354058 47574 354294
rect 46954 320614 47574 354058
rect 46954 320378 46986 320614
rect 47222 320378 47306 320614
rect 47542 320378 47574 320614
rect 46954 320294 47574 320378
rect 46954 320058 46986 320294
rect 47222 320058 47306 320294
rect 47542 320058 47574 320294
rect 46954 286614 47574 320058
rect 46954 286378 46986 286614
rect 47222 286378 47306 286614
rect 47542 286378 47574 286614
rect 46954 286294 47574 286378
rect 46954 286058 46986 286294
rect 47222 286058 47306 286294
rect 47542 286058 47574 286294
rect 46954 252614 47574 286058
rect 46954 252378 46986 252614
rect 47222 252378 47306 252614
rect 47542 252378 47574 252614
rect 46954 252294 47574 252378
rect 46954 252058 46986 252294
rect 47222 252058 47306 252294
rect 47542 252058 47574 252294
rect 46954 225560 47574 252058
rect 50674 708678 51294 711590
rect 50674 708442 50706 708678
rect 50942 708442 51026 708678
rect 51262 708442 51294 708678
rect 50674 708358 51294 708442
rect 50674 708122 50706 708358
rect 50942 708122 51026 708358
rect 51262 708122 51294 708358
rect 50674 698334 51294 708122
rect 50674 698098 50706 698334
rect 50942 698098 51026 698334
rect 51262 698098 51294 698334
rect 50674 698014 51294 698098
rect 50674 697778 50706 698014
rect 50942 697778 51026 698014
rect 51262 697778 51294 698014
rect 50674 664334 51294 697778
rect 50674 664098 50706 664334
rect 50942 664098 51026 664334
rect 51262 664098 51294 664334
rect 50674 664014 51294 664098
rect 50674 663778 50706 664014
rect 50942 663778 51026 664014
rect 51262 663778 51294 664014
rect 50674 630334 51294 663778
rect 50674 630098 50706 630334
rect 50942 630098 51026 630334
rect 51262 630098 51294 630334
rect 50674 630014 51294 630098
rect 50674 629778 50706 630014
rect 50942 629778 51026 630014
rect 51262 629778 51294 630014
rect 50674 596334 51294 629778
rect 50674 596098 50706 596334
rect 50942 596098 51026 596334
rect 51262 596098 51294 596334
rect 50674 596014 51294 596098
rect 50674 595778 50706 596014
rect 50942 595778 51026 596014
rect 51262 595778 51294 596014
rect 50674 562334 51294 595778
rect 50674 562098 50706 562334
rect 50942 562098 51026 562334
rect 51262 562098 51294 562334
rect 50674 562014 51294 562098
rect 50674 561778 50706 562014
rect 50942 561778 51026 562014
rect 51262 561778 51294 562014
rect 50674 528334 51294 561778
rect 50674 528098 50706 528334
rect 50942 528098 51026 528334
rect 51262 528098 51294 528334
rect 50674 528014 51294 528098
rect 50674 527778 50706 528014
rect 50942 527778 51026 528014
rect 51262 527778 51294 528014
rect 50674 494334 51294 527778
rect 50674 494098 50706 494334
rect 50942 494098 51026 494334
rect 51262 494098 51294 494334
rect 50674 494014 51294 494098
rect 50674 493778 50706 494014
rect 50942 493778 51026 494014
rect 51262 493778 51294 494014
rect 50674 460334 51294 493778
rect 50674 460098 50706 460334
rect 50942 460098 51026 460334
rect 51262 460098 51294 460334
rect 50674 460014 51294 460098
rect 50674 459778 50706 460014
rect 50942 459778 51026 460014
rect 51262 459778 51294 460014
rect 50674 426334 51294 459778
rect 50674 426098 50706 426334
rect 50942 426098 51026 426334
rect 51262 426098 51294 426334
rect 50674 426014 51294 426098
rect 50674 425778 50706 426014
rect 50942 425778 51026 426014
rect 51262 425778 51294 426014
rect 50674 392334 51294 425778
rect 50674 392098 50706 392334
rect 50942 392098 51026 392334
rect 51262 392098 51294 392334
rect 50674 392014 51294 392098
rect 50674 391778 50706 392014
rect 50942 391778 51026 392014
rect 51262 391778 51294 392014
rect 50674 358334 51294 391778
rect 50674 358098 50706 358334
rect 50942 358098 51026 358334
rect 51262 358098 51294 358334
rect 50674 358014 51294 358098
rect 50674 357778 50706 358014
rect 50942 357778 51026 358014
rect 51262 357778 51294 358014
rect 50674 324334 51294 357778
rect 50674 324098 50706 324334
rect 50942 324098 51026 324334
rect 51262 324098 51294 324334
rect 50674 324014 51294 324098
rect 50674 323778 50706 324014
rect 50942 323778 51026 324014
rect 51262 323778 51294 324014
rect 50674 290334 51294 323778
rect 50674 290098 50706 290334
rect 50942 290098 51026 290334
rect 51262 290098 51294 290334
rect 50674 290014 51294 290098
rect 50674 289778 50706 290014
rect 50942 289778 51026 290014
rect 51262 289778 51294 290014
rect 50674 256334 51294 289778
rect 50674 256098 50706 256334
rect 50942 256098 51026 256334
rect 51262 256098 51294 256334
rect 50674 256014 51294 256098
rect 50674 255778 50706 256014
rect 50942 255778 51026 256014
rect 51262 255778 51294 256014
rect 50674 225560 51294 255778
rect 54394 709638 55014 711590
rect 54394 709402 54426 709638
rect 54662 709402 54746 709638
rect 54982 709402 55014 709638
rect 54394 709318 55014 709402
rect 54394 709082 54426 709318
rect 54662 709082 54746 709318
rect 54982 709082 55014 709318
rect 54394 668054 55014 709082
rect 54394 667818 54426 668054
rect 54662 667818 54746 668054
rect 54982 667818 55014 668054
rect 54394 667734 55014 667818
rect 54394 667498 54426 667734
rect 54662 667498 54746 667734
rect 54982 667498 55014 667734
rect 54394 634054 55014 667498
rect 54394 633818 54426 634054
rect 54662 633818 54746 634054
rect 54982 633818 55014 634054
rect 54394 633734 55014 633818
rect 54394 633498 54426 633734
rect 54662 633498 54746 633734
rect 54982 633498 55014 633734
rect 54394 600054 55014 633498
rect 54394 599818 54426 600054
rect 54662 599818 54746 600054
rect 54982 599818 55014 600054
rect 54394 599734 55014 599818
rect 54394 599498 54426 599734
rect 54662 599498 54746 599734
rect 54982 599498 55014 599734
rect 54394 566054 55014 599498
rect 54394 565818 54426 566054
rect 54662 565818 54746 566054
rect 54982 565818 55014 566054
rect 54394 565734 55014 565818
rect 54394 565498 54426 565734
rect 54662 565498 54746 565734
rect 54982 565498 55014 565734
rect 54394 532054 55014 565498
rect 54394 531818 54426 532054
rect 54662 531818 54746 532054
rect 54982 531818 55014 532054
rect 54394 531734 55014 531818
rect 54394 531498 54426 531734
rect 54662 531498 54746 531734
rect 54982 531498 55014 531734
rect 54394 498054 55014 531498
rect 54394 497818 54426 498054
rect 54662 497818 54746 498054
rect 54982 497818 55014 498054
rect 54394 497734 55014 497818
rect 54394 497498 54426 497734
rect 54662 497498 54746 497734
rect 54982 497498 55014 497734
rect 54394 464054 55014 497498
rect 54394 463818 54426 464054
rect 54662 463818 54746 464054
rect 54982 463818 55014 464054
rect 54394 463734 55014 463818
rect 54394 463498 54426 463734
rect 54662 463498 54746 463734
rect 54982 463498 55014 463734
rect 54394 430054 55014 463498
rect 54394 429818 54426 430054
rect 54662 429818 54746 430054
rect 54982 429818 55014 430054
rect 54394 429734 55014 429818
rect 54394 429498 54426 429734
rect 54662 429498 54746 429734
rect 54982 429498 55014 429734
rect 54394 396054 55014 429498
rect 54394 395818 54426 396054
rect 54662 395818 54746 396054
rect 54982 395818 55014 396054
rect 54394 395734 55014 395818
rect 54394 395498 54426 395734
rect 54662 395498 54746 395734
rect 54982 395498 55014 395734
rect 54394 362054 55014 395498
rect 54394 361818 54426 362054
rect 54662 361818 54746 362054
rect 54982 361818 55014 362054
rect 54394 361734 55014 361818
rect 54394 361498 54426 361734
rect 54662 361498 54746 361734
rect 54982 361498 55014 361734
rect 54394 328054 55014 361498
rect 54394 327818 54426 328054
rect 54662 327818 54746 328054
rect 54982 327818 55014 328054
rect 54394 327734 55014 327818
rect 54394 327498 54426 327734
rect 54662 327498 54746 327734
rect 54982 327498 55014 327734
rect 54394 294054 55014 327498
rect 54394 293818 54426 294054
rect 54662 293818 54746 294054
rect 54982 293818 55014 294054
rect 54394 293734 55014 293818
rect 54394 293498 54426 293734
rect 54662 293498 54746 293734
rect 54982 293498 55014 293734
rect 54394 260054 55014 293498
rect 54394 259818 54426 260054
rect 54662 259818 54746 260054
rect 54982 259818 55014 260054
rect 54394 259734 55014 259818
rect 54394 259498 54426 259734
rect 54662 259498 54746 259734
rect 54982 259498 55014 259734
rect 54394 225941 55014 259498
rect 54394 225705 54426 225941
rect 54662 225705 54746 225941
rect 54982 225705 55014 225941
rect 54394 225560 55014 225705
rect 58114 710598 58734 711590
rect 58114 710362 58146 710598
rect 58382 710362 58466 710598
rect 58702 710362 58734 710598
rect 58114 710278 58734 710362
rect 58114 710042 58146 710278
rect 58382 710042 58466 710278
rect 58702 710042 58734 710278
rect 58114 671774 58734 710042
rect 58114 671538 58146 671774
rect 58382 671538 58466 671774
rect 58702 671538 58734 671774
rect 58114 671454 58734 671538
rect 58114 671218 58146 671454
rect 58382 671218 58466 671454
rect 58702 671218 58734 671454
rect 58114 637774 58734 671218
rect 58114 637538 58146 637774
rect 58382 637538 58466 637774
rect 58702 637538 58734 637774
rect 58114 637454 58734 637538
rect 58114 637218 58146 637454
rect 58382 637218 58466 637454
rect 58702 637218 58734 637454
rect 58114 603774 58734 637218
rect 58114 603538 58146 603774
rect 58382 603538 58466 603774
rect 58702 603538 58734 603774
rect 58114 603454 58734 603538
rect 58114 603218 58146 603454
rect 58382 603218 58466 603454
rect 58702 603218 58734 603454
rect 58114 569774 58734 603218
rect 58114 569538 58146 569774
rect 58382 569538 58466 569774
rect 58702 569538 58734 569774
rect 58114 569454 58734 569538
rect 58114 569218 58146 569454
rect 58382 569218 58466 569454
rect 58702 569218 58734 569454
rect 58114 535774 58734 569218
rect 58114 535538 58146 535774
rect 58382 535538 58466 535774
rect 58702 535538 58734 535774
rect 58114 535454 58734 535538
rect 58114 535218 58146 535454
rect 58382 535218 58466 535454
rect 58702 535218 58734 535454
rect 58114 501774 58734 535218
rect 58114 501538 58146 501774
rect 58382 501538 58466 501774
rect 58702 501538 58734 501774
rect 58114 501454 58734 501538
rect 58114 501218 58146 501454
rect 58382 501218 58466 501454
rect 58702 501218 58734 501454
rect 58114 467774 58734 501218
rect 58114 467538 58146 467774
rect 58382 467538 58466 467774
rect 58702 467538 58734 467774
rect 58114 467454 58734 467538
rect 58114 467218 58146 467454
rect 58382 467218 58466 467454
rect 58702 467218 58734 467454
rect 58114 433774 58734 467218
rect 58114 433538 58146 433774
rect 58382 433538 58466 433774
rect 58702 433538 58734 433774
rect 58114 433454 58734 433538
rect 58114 433218 58146 433454
rect 58382 433218 58466 433454
rect 58702 433218 58734 433454
rect 58114 399774 58734 433218
rect 58114 399538 58146 399774
rect 58382 399538 58466 399774
rect 58702 399538 58734 399774
rect 58114 399454 58734 399538
rect 58114 399218 58146 399454
rect 58382 399218 58466 399454
rect 58702 399218 58734 399454
rect 58114 365774 58734 399218
rect 58114 365538 58146 365774
rect 58382 365538 58466 365774
rect 58702 365538 58734 365774
rect 58114 365454 58734 365538
rect 58114 365218 58146 365454
rect 58382 365218 58466 365454
rect 58702 365218 58734 365454
rect 58114 331774 58734 365218
rect 58114 331538 58146 331774
rect 58382 331538 58466 331774
rect 58702 331538 58734 331774
rect 58114 331454 58734 331538
rect 58114 331218 58146 331454
rect 58382 331218 58466 331454
rect 58702 331218 58734 331454
rect 58114 297774 58734 331218
rect 58114 297538 58146 297774
rect 58382 297538 58466 297774
rect 58702 297538 58734 297774
rect 58114 297454 58734 297538
rect 58114 297218 58146 297454
rect 58382 297218 58466 297454
rect 58702 297218 58734 297454
rect 58114 263774 58734 297218
rect 58114 263538 58146 263774
rect 58382 263538 58466 263774
rect 58702 263538 58734 263774
rect 58114 263454 58734 263538
rect 58114 263218 58146 263454
rect 58382 263218 58466 263454
rect 58702 263218 58734 263454
rect 58114 229774 58734 263218
rect 58114 229538 58146 229774
rect 58382 229538 58466 229774
rect 58702 229538 58734 229774
rect 58114 229454 58734 229538
rect 58114 229218 58146 229454
rect 58382 229218 58466 229454
rect 58702 229218 58734 229454
rect 58114 225560 58734 229218
rect 61834 711558 62454 711590
rect 61834 711322 61866 711558
rect 62102 711322 62186 711558
rect 62422 711322 62454 711558
rect 61834 711238 62454 711322
rect 61834 711002 61866 711238
rect 62102 711002 62186 711238
rect 62422 711002 62454 711238
rect 61834 675494 62454 711002
rect 61834 675258 61866 675494
rect 62102 675258 62186 675494
rect 62422 675258 62454 675494
rect 61834 675174 62454 675258
rect 61834 674938 61866 675174
rect 62102 674938 62186 675174
rect 62422 674938 62454 675174
rect 61834 641494 62454 674938
rect 61834 641258 61866 641494
rect 62102 641258 62186 641494
rect 62422 641258 62454 641494
rect 61834 641174 62454 641258
rect 61834 640938 61866 641174
rect 62102 640938 62186 641174
rect 62422 640938 62454 641174
rect 61834 607494 62454 640938
rect 61834 607258 61866 607494
rect 62102 607258 62186 607494
rect 62422 607258 62454 607494
rect 61834 607174 62454 607258
rect 61834 606938 61866 607174
rect 62102 606938 62186 607174
rect 62422 606938 62454 607174
rect 61834 573494 62454 606938
rect 61834 573258 61866 573494
rect 62102 573258 62186 573494
rect 62422 573258 62454 573494
rect 61834 573174 62454 573258
rect 61834 572938 61866 573174
rect 62102 572938 62186 573174
rect 62422 572938 62454 573174
rect 61834 539494 62454 572938
rect 61834 539258 61866 539494
rect 62102 539258 62186 539494
rect 62422 539258 62454 539494
rect 61834 539174 62454 539258
rect 61834 538938 61866 539174
rect 62102 538938 62186 539174
rect 62422 538938 62454 539174
rect 61834 505494 62454 538938
rect 61834 505258 61866 505494
rect 62102 505258 62186 505494
rect 62422 505258 62454 505494
rect 61834 505174 62454 505258
rect 61834 504938 61866 505174
rect 62102 504938 62186 505174
rect 62422 504938 62454 505174
rect 61834 471494 62454 504938
rect 61834 471258 61866 471494
rect 62102 471258 62186 471494
rect 62422 471258 62454 471494
rect 61834 471174 62454 471258
rect 61834 470938 61866 471174
rect 62102 470938 62186 471174
rect 62422 470938 62454 471174
rect 61834 437494 62454 470938
rect 61834 437258 61866 437494
rect 62102 437258 62186 437494
rect 62422 437258 62454 437494
rect 61834 437174 62454 437258
rect 61834 436938 61866 437174
rect 62102 436938 62186 437174
rect 62422 436938 62454 437174
rect 61834 403494 62454 436938
rect 61834 403258 61866 403494
rect 62102 403258 62186 403494
rect 62422 403258 62454 403494
rect 61834 403174 62454 403258
rect 61834 402938 61866 403174
rect 62102 402938 62186 403174
rect 62422 402938 62454 403174
rect 61834 369494 62454 402938
rect 61834 369258 61866 369494
rect 62102 369258 62186 369494
rect 62422 369258 62454 369494
rect 61834 369174 62454 369258
rect 61834 368938 61866 369174
rect 62102 368938 62186 369174
rect 62422 368938 62454 369174
rect 61834 335494 62454 368938
rect 61834 335258 61866 335494
rect 62102 335258 62186 335494
rect 62422 335258 62454 335494
rect 61834 335174 62454 335258
rect 61834 334938 61866 335174
rect 62102 334938 62186 335174
rect 62422 334938 62454 335174
rect 61834 301494 62454 334938
rect 61834 301258 61866 301494
rect 62102 301258 62186 301494
rect 62422 301258 62454 301494
rect 61834 301174 62454 301258
rect 61834 300938 61866 301174
rect 62102 300938 62186 301174
rect 62422 300938 62454 301174
rect 61834 267494 62454 300938
rect 61834 267258 61866 267494
rect 62102 267258 62186 267494
rect 62422 267258 62454 267494
rect 61834 267174 62454 267258
rect 61834 266938 61866 267174
rect 62102 266938 62186 267174
rect 62422 266938 62454 267174
rect 61834 233494 62454 266938
rect 61834 233258 61866 233494
rect 62102 233258 62186 233494
rect 62422 233258 62454 233494
rect 61834 233174 62454 233258
rect 61834 232938 61866 233174
rect 62102 232938 62186 233174
rect 62422 232938 62454 233174
rect 61834 225560 62454 232938
rect 69794 704838 70414 711590
rect 69794 704602 69826 704838
rect 70062 704602 70146 704838
rect 70382 704602 70414 704838
rect 69794 704518 70414 704602
rect 69794 704282 69826 704518
rect 70062 704282 70146 704518
rect 70382 704282 70414 704518
rect 69794 683454 70414 704282
rect 69794 683218 69826 683454
rect 70062 683218 70146 683454
rect 70382 683218 70414 683454
rect 69794 683134 70414 683218
rect 69794 682898 69826 683134
rect 70062 682898 70146 683134
rect 70382 682898 70414 683134
rect 69794 649454 70414 682898
rect 69794 649218 69826 649454
rect 70062 649218 70146 649454
rect 70382 649218 70414 649454
rect 69794 649134 70414 649218
rect 69794 648898 69826 649134
rect 70062 648898 70146 649134
rect 70382 648898 70414 649134
rect 69794 615454 70414 648898
rect 69794 615218 69826 615454
rect 70062 615218 70146 615454
rect 70382 615218 70414 615454
rect 69794 615134 70414 615218
rect 69794 614898 69826 615134
rect 70062 614898 70146 615134
rect 70382 614898 70414 615134
rect 69794 581454 70414 614898
rect 69794 581218 69826 581454
rect 70062 581218 70146 581454
rect 70382 581218 70414 581454
rect 69794 581134 70414 581218
rect 69794 580898 69826 581134
rect 70062 580898 70146 581134
rect 70382 580898 70414 581134
rect 69794 547454 70414 580898
rect 69794 547218 69826 547454
rect 70062 547218 70146 547454
rect 70382 547218 70414 547454
rect 69794 547134 70414 547218
rect 69794 546898 69826 547134
rect 70062 546898 70146 547134
rect 70382 546898 70414 547134
rect 69794 513454 70414 546898
rect 69794 513218 69826 513454
rect 70062 513218 70146 513454
rect 70382 513218 70414 513454
rect 69794 513134 70414 513218
rect 69794 512898 69826 513134
rect 70062 512898 70146 513134
rect 70382 512898 70414 513134
rect 69794 479454 70414 512898
rect 69794 479218 69826 479454
rect 70062 479218 70146 479454
rect 70382 479218 70414 479454
rect 69794 479134 70414 479218
rect 69794 478898 69826 479134
rect 70062 478898 70146 479134
rect 70382 478898 70414 479134
rect 69794 445454 70414 478898
rect 69794 445218 69826 445454
rect 70062 445218 70146 445454
rect 70382 445218 70414 445454
rect 69794 445134 70414 445218
rect 69794 444898 69826 445134
rect 70062 444898 70146 445134
rect 70382 444898 70414 445134
rect 69794 411454 70414 444898
rect 69794 411218 69826 411454
rect 70062 411218 70146 411454
rect 70382 411218 70414 411454
rect 69794 411134 70414 411218
rect 69794 410898 69826 411134
rect 70062 410898 70146 411134
rect 70382 410898 70414 411134
rect 69794 377454 70414 410898
rect 69794 377218 69826 377454
rect 70062 377218 70146 377454
rect 70382 377218 70414 377454
rect 69794 377134 70414 377218
rect 69794 376898 69826 377134
rect 70062 376898 70146 377134
rect 70382 376898 70414 377134
rect 69794 343454 70414 376898
rect 69794 343218 69826 343454
rect 70062 343218 70146 343454
rect 70382 343218 70414 343454
rect 69794 343134 70414 343218
rect 69794 342898 69826 343134
rect 70062 342898 70146 343134
rect 70382 342898 70414 343134
rect 69794 309454 70414 342898
rect 69794 309218 69826 309454
rect 70062 309218 70146 309454
rect 70382 309218 70414 309454
rect 69794 309134 70414 309218
rect 69794 308898 69826 309134
rect 70062 308898 70146 309134
rect 70382 308898 70414 309134
rect 69794 275454 70414 308898
rect 69794 275218 69826 275454
rect 70062 275218 70146 275454
rect 70382 275218 70414 275454
rect 69794 275134 70414 275218
rect 69794 274898 69826 275134
rect 70062 274898 70146 275134
rect 70382 274898 70414 275134
rect 69794 241454 70414 274898
rect 69794 241218 69826 241454
rect 70062 241218 70146 241454
rect 70382 241218 70414 241454
rect 69794 241134 70414 241218
rect 69794 240898 69826 241134
rect 70062 240898 70146 241134
rect 70382 240898 70414 241134
rect 69794 232680 70414 240898
rect 73514 705798 74134 711590
rect 73514 705562 73546 705798
rect 73782 705562 73866 705798
rect 74102 705562 74134 705798
rect 73514 705478 74134 705562
rect 73514 705242 73546 705478
rect 73782 705242 73866 705478
rect 74102 705242 74134 705478
rect 73514 687174 74134 705242
rect 73514 686938 73546 687174
rect 73782 686938 73866 687174
rect 74102 686938 74134 687174
rect 73514 686854 74134 686938
rect 73514 686618 73546 686854
rect 73782 686618 73866 686854
rect 74102 686618 74134 686854
rect 73514 653174 74134 686618
rect 73514 652938 73546 653174
rect 73782 652938 73866 653174
rect 74102 652938 74134 653174
rect 73514 652854 74134 652938
rect 73514 652618 73546 652854
rect 73782 652618 73866 652854
rect 74102 652618 74134 652854
rect 73514 619174 74134 652618
rect 73514 618938 73546 619174
rect 73782 618938 73866 619174
rect 74102 618938 74134 619174
rect 73514 618854 74134 618938
rect 73514 618618 73546 618854
rect 73782 618618 73866 618854
rect 74102 618618 74134 618854
rect 73514 585174 74134 618618
rect 73514 584938 73546 585174
rect 73782 584938 73866 585174
rect 74102 584938 74134 585174
rect 73514 584854 74134 584938
rect 73514 584618 73546 584854
rect 73782 584618 73866 584854
rect 74102 584618 74134 584854
rect 73514 551174 74134 584618
rect 73514 550938 73546 551174
rect 73782 550938 73866 551174
rect 74102 550938 74134 551174
rect 73514 550854 74134 550938
rect 73514 550618 73546 550854
rect 73782 550618 73866 550854
rect 74102 550618 74134 550854
rect 73514 517174 74134 550618
rect 73514 516938 73546 517174
rect 73782 516938 73866 517174
rect 74102 516938 74134 517174
rect 73514 516854 74134 516938
rect 73514 516618 73546 516854
rect 73782 516618 73866 516854
rect 74102 516618 74134 516854
rect 73514 483174 74134 516618
rect 73514 482938 73546 483174
rect 73782 482938 73866 483174
rect 74102 482938 74134 483174
rect 73514 482854 74134 482938
rect 73514 482618 73546 482854
rect 73782 482618 73866 482854
rect 74102 482618 74134 482854
rect 73514 449174 74134 482618
rect 73514 448938 73546 449174
rect 73782 448938 73866 449174
rect 74102 448938 74134 449174
rect 73514 448854 74134 448938
rect 73514 448618 73546 448854
rect 73782 448618 73866 448854
rect 74102 448618 74134 448854
rect 73514 415174 74134 448618
rect 73514 414938 73546 415174
rect 73782 414938 73866 415174
rect 74102 414938 74134 415174
rect 73514 414854 74134 414938
rect 73514 414618 73546 414854
rect 73782 414618 73866 414854
rect 74102 414618 74134 414854
rect 73514 381174 74134 414618
rect 73514 380938 73546 381174
rect 73782 380938 73866 381174
rect 74102 380938 74134 381174
rect 73514 380854 74134 380938
rect 73514 380618 73546 380854
rect 73782 380618 73866 380854
rect 74102 380618 74134 380854
rect 73514 347174 74134 380618
rect 73514 346938 73546 347174
rect 73782 346938 73866 347174
rect 74102 346938 74134 347174
rect 73514 346854 74134 346938
rect 73514 346618 73546 346854
rect 73782 346618 73866 346854
rect 74102 346618 74134 346854
rect 73514 313174 74134 346618
rect 73514 312938 73546 313174
rect 73782 312938 73866 313174
rect 74102 312938 74134 313174
rect 73514 312854 74134 312938
rect 73514 312618 73546 312854
rect 73782 312618 73866 312854
rect 74102 312618 74134 312854
rect 73514 279174 74134 312618
rect 73514 278938 73546 279174
rect 73782 278938 73866 279174
rect 74102 278938 74134 279174
rect 73514 278854 74134 278938
rect 73514 278618 73546 278854
rect 73782 278618 73866 278854
rect 74102 278618 74134 278854
rect 73514 245174 74134 278618
rect 73514 244938 73546 245174
rect 73782 244938 73866 245174
rect 74102 244938 74134 245174
rect 73514 244854 74134 244938
rect 73514 244618 73546 244854
rect 73782 244618 73866 244854
rect 74102 244618 74134 244854
rect 65300 229771 70094 229800
rect 65300 229535 65339 229771
rect 65575 229535 65659 229771
rect 65895 229535 65979 229771
rect 66215 229535 66299 229771
rect 66535 229535 66619 229771
rect 66855 229535 66939 229771
rect 67175 229535 67259 229771
rect 67495 229535 67579 229771
rect 67815 229535 67899 229771
rect 68135 229535 68219 229771
rect 68455 229535 68539 229771
rect 68775 229535 68859 229771
rect 69095 229535 69179 229771
rect 69415 229535 69499 229771
rect 69735 229535 69819 229771
rect 70055 229535 70094 229771
rect 65300 229451 70094 229535
rect 65300 229215 65339 229451
rect 65575 229215 65659 229451
rect 65895 229215 65979 229451
rect 66215 229215 66299 229451
rect 66535 229215 66619 229451
rect 66855 229215 66939 229451
rect 67175 229215 67259 229451
rect 67495 229215 67579 229451
rect 67815 229215 67899 229451
rect 68135 229215 68219 229451
rect 68455 229215 68539 229451
rect 68775 229215 68859 229451
rect 69095 229215 69179 229451
rect 69415 229215 69499 229451
rect 69735 229215 69819 229451
rect 70055 229215 70094 229451
rect 65300 229186 70094 229215
rect 65300 225801 71300 225900
rect 65300 225565 65462 225801
rect 65698 225565 65782 225801
rect 66018 225565 66102 225801
rect 66338 225565 66422 225801
rect 66658 225565 66742 225801
rect 66978 225565 67062 225801
rect 67298 225565 67382 225801
rect 67618 225565 67702 225801
rect 67938 225565 68022 225801
rect 68258 225565 68342 225801
rect 68578 225565 68662 225801
rect 68898 225565 68982 225801
rect 69218 225565 69302 225801
rect 69538 225565 69622 225801
rect 69858 225565 69942 225801
rect 70178 225565 70262 225801
rect 70498 225565 70582 225801
rect 70818 225565 70902 225801
rect 71138 225565 71300 225801
rect 73514 225660 74134 244618
rect 77234 706758 77854 711590
rect 77234 706522 77266 706758
rect 77502 706522 77586 706758
rect 77822 706522 77854 706758
rect 77234 706438 77854 706522
rect 77234 706202 77266 706438
rect 77502 706202 77586 706438
rect 77822 706202 77854 706438
rect 77234 690894 77854 706202
rect 77234 690658 77266 690894
rect 77502 690658 77586 690894
rect 77822 690658 77854 690894
rect 77234 690574 77854 690658
rect 77234 690338 77266 690574
rect 77502 690338 77586 690574
rect 77822 690338 77854 690574
rect 77234 656894 77854 690338
rect 77234 656658 77266 656894
rect 77502 656658 77586 656894
rect 77822 656658 77854 656894
rect 77234 656574 77854 656658
rect 77234 656338 77266 656574
rect 77502 656338 77586 656574
rect 77822 656338 77854 656574
rect 77234 622894 77854 656338
rect 77234 622658 77266 622894
rect 77502 622658 77586 622894
rect 77822 622658 77854 622894
rect 77234 622574 77854 622658
rect 77234 622338 77266 622574
rect 77502 622338 77586 622574
rect 77822 622338 77854 622574
rect 77234 588894 77854 622338
rect 77234 588658 77266 588894
rect 77502 588658 77586 588894
rect 77822 588658 77854 588894
rect 77234 588574 77854 588658
rect 77234 588338 77266 588574
rect 77502 588338 77586 588574
rect 77822 588338 77854 588574
rect 77234 554894 77854 588338
rect 77234 554658 77266 554894
rect 77502 554658 77586 554894
rect 77822 554658 77854 554894
rect 77234 554574 77854 554658
rect 77234 554338 77266 554574
rect 77502 554338 77586 554574
rect 77822 554338 77854 554574
rect 77234 520894 77854 554338
rect 77234 520658 77266 520894
rect 77502 520658 77586 520894
rect 77822 520658 77854 520894
rect 77234 520574 77854 520658
rect 77234 520338 77266 520574
rect 77502 520338 77586 520574
rect 77822 520338 77854 520574
rect 77234 486894 77854 520338
rect 77234 486658 77266 486894
rect 77502 486658 77586 486894
rect 77822 486658 77854 486894
rect 77234 486574 77854 486658
rect 77234 486338 77266 486574
rect 77502 486338 77586 486574
rect 77822 486338 77854 486574
rect 77234 452894 77854 486338
rect 77234 452658 77266 452894
rect 77502 452658 77586 452894
rect 77822 452658 77854 452894
rect 77234 452574 77854 452658
rect 77234 452338 77266 452574
rect 77502 452338 77586 452574
rect 77822 452338 77854 452574
rect 77234 418894 77854 452338
rect 77234 418658 77266 418894
rect 77502 418658 77586 418894
rect 77822 418658 77854 418894
rect 77234 418574 77854 418658
rect 77234 418338 77266 418574
rect 77502 418338 77586 418574
rect 77822 418338 77854 418574
rect 77234 384894 77854 418338
rect 77234 384658 77266 384894
rect 77502 384658 77586 384894
rect 77822 384658 77854 384894
rect 77234 384574 77854 384658
rect 77234 384338 77266 384574
rect 77502 384338 77586 384574
rect 77822 384338 77854 384574
rect 77234 350894 77854 384338
rect 77234 350658 77266 350894
rect 77502 350658 77586 350894
rect 77822 350658 77854 350894
rect 77234 350574 77854 350658
rect 77234 350338 77266 350574
rect 77502 350338 77586 350574
rect 77822 350338 77854 350574
rect 77234 316894 77854 350338
rect 77234 316658 77266 316894
rect 77502 316658 77586 316894
rect 77822 316658 77854 316894
rect 77234 316574 77854 316658
rect 77234 316338 77266 316574
rect 77502 316338 77586 316574
rect 77822 316338 77854 316574
rect 77234 282894 77854 316338
rect 77234 282658 77266 282894
rect 77502 282658 77586 282894
rect 77822 282658 77854 282894
rect 77234 282574 77854 282658
rect 77234 282338 77266 282574
rect 77502 282338 77586 282574
rect 77822 282338 77854 282574
rect 77234 248894 77854 282338
rect 77234 248658 77266 248894
rect 77502 248658 77586 248894
rect 77822 248658 77854 248894
rect 77234 248574 77854 248658
rect 77234 248338 77266 248574
rect 77502 248338 77586 248574
rect 77822 248338 77854 248574
rect 77234 225660 77854 248338
rect 80954 707718 81574 711590
rect 80954 707482 80986 707718
rect 81222 707482 81306 707718
rect 81542 707482 81574 707718
rect 80954 707398 81574 707482
rect 80954 707162 80986 707398
rect 81222 707162 81306 707398
rect 81542 707162 81574 707398
rect 80954 694614 81574 707162
rect 80954 694378 80986 694614
rect 81222 694378 81306 694614
rect 81542 694378 81574 694614
rect 80954 694294 81574 694378
rect 80954 694058 80986 694294
rect 81222 694058 81306 694294
rect 81542 694058 81574 694294
rect 80954 660614 81574 694058
rect 80954 660378 80986 660614
rect 81222 660378 81306 660614
rect 81542 660378 81574 660614
rect 80954 660294 81574 660378
rect 80954 660058 80986 660294
rect 81222 660058 81306 660294
rect 81542 660058 81574 660294
rect 80954 626614 81574 660058
rect 80954 626378 80986 626614
rect 81222 626378 81306 626614
rect 81542 626378 81574 626614
rect 80954 626294 81574 626378
rect 80954 626058 80986 626294
rect 81222 626058 81306 626294
rect 81542 626058 81574 626294
rect 80954 592614 81574 626058
rect 80954 592378 80986 592614
rect 81222 592378 81306 592614
rect 81542 592378 81574 592614
rect 80954 592294 81574 592378
rect 80954 592058 80986 592294
rect 81222 592058 81306 592294
rect 81542 592058 81574 592294
rect 80954 558614 81574 592058
rect 80954 558378 80986 558614
rect 81222 558378 81306 558614
rect 81542 558378 81574 558614
rect 80954 558294 81574 558378
rect 80954 558058 80986 558294
rect 81222 558058 81306 558294
rect 81542 558058 81574 558294
rect 80954 524614 81574 558058
rect 80954 524378 80986 524614
rect 81222 524378 81306 524614
rect 81542 524378 81574 524614
rect 80954 524294 81574 524378
rect 80954 524058 80986 524294
rect 81222 524058 81306 524294
rect 81542 524058 81574 524294
rect 80954 490614 81574 524058
rect 80954 490378 80986 490614
rect 81222 490378 81306 490614
rect 81542 490378 81574 490614
rect 80954 490294 81574 490378
rect 80954 490058 80986 490294
rect 81222 490058 81306 490294
rect 81542 490058 81574 490294
rect 80954 456614 81574 490058
rect 80954 456378 80986 456614
rect 81222 456378 81306 456614
rect 81542 456378 81574 456614
rect 80954 456294 81574 456378
rect 80954 456058 80986 456294
rect 81222 456058 81306 456294
rect 81542 456058 81574 456294
rect 80954 422614 81574 456058
rect 80954 422378 80986 422614
rect 81222 422378 81306 422614
rect 81542 422378 81574 422614
rect 80954 422294 81574 422378
rect 80954 422058 80986 422294
rect 81222 422058 81306 422294
rect 81542 422058 81574 422294
rect 80954 388614 81574 422058
rect 80954 388378 80986 388614
rect 81222 388378 81306 388614
rect 81542 388378 81574 388614
rect 80954 388294 81574 388378
rect 80954 388058 80986 388294
rect 81222 388058 81306 388294
rect 81542 388058 81574 388294
rect 80954 354614 81574 388058
rect 80954 354378 80986 354614
rect 81222 354378 81306 354614
rect 81542 354378 81574 354614
rect 80954 354294 81574 354378
rect 80954 354058 80986 354294
rect 81222 354058 81306 354294
rect 81542 354058 81574 354294
rect 80954 320614 81574 354058
rect 80954 320378 80986 320614
rect 81222 320378 81306 320614
rect 81542 320378 81574 320614
rect 80954 320294 81574 320378
rect 80954 320058 80986 320294
rect 81222 320058 81306 320294
rect 81542 320058 81574 320294
rect 80954 286614 81574 320058
rect 80954 286378 80986 286614
rect 81222 286378 81306 286614
rect 81542 286378 81574 286614
rect 80954 286294 81574 286378
rect 80954 286058 80986 286294
rect 81222 286058 81306 286294
rect 81542 286058 81574 286294
rect 80954 252614 81574 286058
rect 80954 252378 80986 252614
rect 81222 252378 81306 252614
rect 81542 252378 81574 252614
rect 80954 252294 81574 252378
rect 80954 252058 80986 252294
rect 81222 252058 81306 252294
rect 81542 252058 81574 252294
rect 80954 225660 81574 252058
rect 84674 708678 85294 711590
rect 84674 708442 84706 708678
rect 84942 708442 85026 708678
rect 85262 708442 85294 708678
rect 84674 708358 85294 708442
rect 84674 708122 84706 708358
rect 84942 708122 85026 708358
rect 85262 708122 85294 708358
rect 84674 698334 85294 708122
rect 84674 698098 84706 698334
rect 84942 698098 85026 698334
rect 85262 698098 85294 698334
rect 84674 698014 85294 698098
rect 84674 697778 84706 698014
rect 84942 697778 85026 698014
rect 85262 697778 85294 698014
rect 84674 664334 85294 697778
rect 84674 664098 84706 664334
rect 84942 664098 85026 664334
rect 85262 664098 85294 664334
rect 84674 664014 85294 664098
rect 84674 663778 84706 664014
rect 84942 663778 85026 664014
rect 85262 663778 85294 664014
rect 84674 630334 85294 663778
rect 84674 630098 84706 630334
rect 84942 630098 85026 630334
rect 85262 630098 85294 630334
rect 84674 630014 85294 630098
rect 84674 629778 84706 630014
rect 84942 629778 85026 630014
rect 85262 629778 85294 630014
rect 84674 596334 85294 629778
rect 84674 596098 84706 596334
rect 84942 596098 85026 596334
rect 85262 596098 85294 596334
rect 84674 596014 85294 596098
rect 84674 595778 84706 596014
rect 84942 595778 85026 596014
rect 85262 595778 85294 596014
rect 84674 562334 85294 595778
rect 84674 562098 84706 562334
rect 84942 562098 85026 562334
rect 85262 562098 85294 562334
rect 84674 562014 85294 562098
rect 84674 561778 84706 562014
rect 84942 561778 85026 562014
rect 85262 561778 85294 562014
rect 84674 528334 85294 561778
rect 84674 528098 84706 528334
rect 84942 528098 85026 528334
rect 85262 528098 85294 528334
rect 84674 528014 85294 528098
rect 84674 527778 84706 528014
rect 84942 527778 85026 528014
rect 85262 527778 85294 528014
rect 84674 494334 85294 527778
rect 84674 494098 84706 494334
rect 84942 494098 85026 494334
rect 85262 494098 85294 494334
rect 84674 494014 85294 494098
rect 84674 493778 84706 494014
rect 84942 493778 85026 494014
rect 85262 493778 85294 494014
rect 84674 460334 85294 493778
rect 84674 460098 84706 460334
rect 84942 460098 85026 460334
rect 85262 460098 85294 460334
rect 84674 460014 85294 460098
rect 84674 459778 84706 460014
rect 84942 459778 85026 460014
rect 85262 459778 85294 460014
rect 84674 426334 85294 459778
rect 84674 426098 84706 426334
rect 84942 426098 85026 426334
rect 85262 426098 85294 426334
rect 84674 426014 85294 426098
rect 84674 425778 84706 426014
rect 84942 425778 85026 426014
rect 85262 425778 85294 426014
rect 84674 392334 85294 425778
rect 84674 392098 84706 392334
rect 84942 392098 85026 392334
rect 85262 392098 85294 392334
rect 84674 392014 85294 392098
rect 84674 391778 84706 392014
rect 84942 391778 85026 392014
rect 85262 391778 85294 392014
rect 84674 358334 85294 391778
rect 84674 358098 84706 358334
rect 84942 358098 85026 358334
rect 85262 358098 85294 358334
rect 84674 358014 85294 358098
rect 84674 357778 84706 358014
rect 84942 357778 85026 358014
rect 85262 357778 85294 358014
rect 84674 324334 85294 357778
rect 84674 324098 84706 324334
rect 84942 324098 85026 324334
rect 85262 324098 85294 324334
rect 84674 324014 85294 324098
rect 84674 323778 84706 324014
rect 84942 323778 85026 324014
rect 85262 323778 85294 324014
rect 84674 290334 85294 323778
rect 84674 290098 84706 290334
rect 84942 290098 85026 290334
rect 85262 290098 85294 290334
rect 84674 290014 85294 290098
rect 84674 289778 84706 290014
rect 84942 289778 85026 290014
rect 85262 289778 85294 290014
rect 84674 256334 85294 289778
rect 84674 256098 84706 256334
rect 84942 256098 85026 256334
rect 85262 256098 85294 256334
rect 84674 256014 85294 256098
rect 84674 255778 84706 256014
rect 84942 255778 85026 256014
rect 85262 255778 85294 256014
rect 84674 225660 85294 255778
rect 88394 709638 89014 711590
rect 88394 709402 88426 709638
rect 88662 709402 88746 709638
rect 88982 709402 89014 709638
rect 88394 709318 89014 709402
rect 88394 709082 88426 709318
rect 88662 709082 88746 709318
rect 88982 709082 89014 709318
rect 88394 668054 89014 709082
rect 88394 667818 88426 668054
rect 88662 667818 88746 668054
rect 88982 667818 89014 668054
rect 88394 667734 89014 667818
rect 88394 667498 88426 667734
rect 88662 667498 88746 667734
rect 88982 667498 89014 667734
rect 88394 634054 89014 667498
rect 88394 633818 88426 634054
rect 88662 633818 88746 634054
rect 88982 633818 89014 634054
rect 88394 633734 89014 633818
rect 88394 633498 88426 633734
rect 88662 633498 88746 633734
rect 88982 633498 89014 633734
rect 88394 600054 89014 633498
rect 88394 599818 88426 600054
rect 88662 599818 88746 600054
rect 88982 599818 89014 600054
rect 88394 599734 89014 599818
rect 88394 599498 88426 599734
rect 88662 599498 88746 599734
rect 88982 599498 89014 599734
rect 88394 566054 89014 599498
rect 88394 565818 88426 566054
rect 88662 565818 88746 566054
rect 88982 565818 89014 566054
rect 88394 565734 89014 565818
rect 88394 565498 88426 565734
rect 88662 565498 88746 565734
rect 88982 565498 89014 565734
rect 88394 532054 89014 565498
rect 88394 531818 88426 532054
rect 88662 531818 88746 532054
rect 88982 531818 89014 532054
rect 88394 531734 89014 531818
rect 88394 531498 88426 531734
rect 88662 531498 88746 531734
rect 88982 531498 89014 531734
rect 88394 498054 89014 531498
rect 88394 497818 88426 498054
rect 88662 497818 88746 498054
rect 88982 497818 89014 498054
rect 88394 497734 89014 497818
rect 88394 497498 88426 497734
rect 88662 497498 88746 497734
rect 88982 497498 89014 497734
rect 88394 464054 89014 497498
rect 88394 463818 88426 464054
rect 88662 463818 88746 464054
rect 88982 463818 89014 464054
rect 88394 463734 89014 463818
rect 88394 463498 88426 463734
rect 88662 463498 88746 463734
rect 88982 463498 89014 463734
rect 88394 430054 89014 463498
rect 88394 429818 88426 430054
rect 88662 429818 88746 430054
rect 88982 429818 89014 430054
rect 88394 429734 89014 429818
rect 88394 429498 88426 429734
rect 88662 429498 88746 429734
rect 88982 429498 89014 429734
rect 88394 396054 89014 429498
rect 88394 395818 88426 396054
rect 88662 395818 88746 396054
rect 88982 395818 89014 396054
rect 88394 395734 89014 395818
rect 88394 395498 88426 395734
rect 88662 395498 88746 395734
rect 88982 395498 89014 395734
rect 88394 362054 89014 395498
rect 88394 361818 88426 362054
rect 88662 361818 88746 362054
rect 88982 361818 89014 362054
rect 88394 361734 89014 361818
rect 88394 361498 88426 361734
rect 88662 361498 88746 361734
rect 88982 361498 89014 361734
rect 88394 328054 89014 361498
rect 88394 327818 88426 328054
rect 88662 327818 88746 328054
rect 88982 327818 89014 328054
rect 88394 327734 89014 327818
rect 88394 327498 88426 327734
rect 88662 327498 88746 327734
rect 88982 327498 89014 327734
rect 88394 294054 89014 327498
rect 88394 293818 88426 294054
rect 88662 293818 88746 294054
rect 88982 293818 89014 294054
rect 88394 293734 89014 293818
rect 88394 293498 88426 293734
rect 88662 293498 88746 293734
rect 88982 293498 89014 293734
rect 88394 260054 89014 293498
rect 88394 259818 88426 260054
rect 88662 259818 88746 260054
rect 88982 259818 89014 260054
rect 88394 259734 89014 259818
rect 88394 259498 88426 259734
rect 88662 259498 88746 259734
rect 88982 259498 89014 259734
rect 88394 225991 89014 259498
rect 88394 225755 88426 225991
rect 88662 225755 88746 225991
rect 88982 225755 89014 225991
rect 88394 225660 89014 225755
rect 92114 710598 92734 711590
rect 92114 710362 92146 710598
rect 92382 710362 92466 710598
rect 92702 710362 92734 710598
rect 92114 710278 92734 710362
rect 92114 710042 92146 710278
rect 92382 710042 92466 710278
rect 92702 710042 92734 710278
rect 92114 671774 92734 710042
rect 92114 671538 92146 671774
rect 92382 671538 92466 671774
rect 92702 671538 92734 671774
rect 92114 671454 92734 671538
rect 92114 671218 92146 671454
rect 92382 671218 92466 671454
rect 92702 671218 92734 671454
rect 92114 637774 92734 671218
rect 92114 637538 92146 637774
rect 92382 637538 92466 637774
rect 92702 637538 92734 637774
rect 92114 637454 92734 637538
rect 92114 637218 92146 637454
rect 92382 637218 92466 637454
rect 92702 637218 92734 637454
rect 92114 603774 92734 637218
rect 92114 603538 92146 603774
rect 92382 603538 92466 603774
rect 92702 603538 92734 603774
rect 92114 603454 92734 603538
rect 92114 603218 92146 603454
rect 92382 603218 92466 603454
rect 92702 603218 92734 603454
rect 92114 569774 92734 603218
rect 92114 569538 92146 569774
rect 92382 569538 92466 569774
rect 92702 569538 92734 569774
rect 92114 569454 92734 569538
rect 92114 569218 92146 569454
rect 92382 569218 92466 569454
rect 92702 569218 92734 569454
rect 92114 535774 92734 569218
rect 92114 535538 92146 535774
rect 92382 535538 92466 535774
rect 92702 535538 92734 535774
rect 92114 535454 92734 535538
rect 92114 535218 92146 535454
rect 92382 535218 92466 535454
rect 92702 535218 92734 535454
rect 92114 501774 92734 535218
rect 92114 501538 92146 501774
rect 92382 501538 92466 501774
rect 92702 501538 92734 501774
rect 92114 501454 92734 501538
rect 92114 501218 92146 501454
rect 92382 501218 92466 501454
rect 92702 501218 92734 501454
rect 92114 467774 92734 501218
rect 92114 467538 92146 467774
rect 92382 467538 92466 467774
rect 92702 467538 92734 467774
rect 92114 467454 92734 467538
rect 92114 467218 92146 467454
rect 92382 467218 92466 467454
rect 92702 467218 92734 467454
rect 92114 433774 92734 467218
rect 92114 433538 92146 433774
rect 92382 433538 92466 433774
rect 92702 433538 92734 433774
rect 92114 433454 92734 433538
rect 92114 433218 92146 433454
rect 92382 433218 92466 433454
rect 92702 433218 92734 433454
rect 92114 399774 92734 433218
rect 92114 399538 92146 399774
rect 92382 399538 92466 399774
rect 92702 399538 92734 399774
rect 92114 399454 92734 399538
rect 92114 399218 92146 399454
rect 92382 399218 92466 399454
rect 92702 399218 92734 399454
rect 92114 365774 92734 399218
rect 92114 365538 92146 365774
rect 92382 365538 92466 365774
rect 92702 365538 92734 365774
rect 92114 365454 92734 365538
rect 92114 365218 92146 365454
rect 92382 365218 92466 365454
rect 92702 365218 92734 365454
rect 92114 331774 92734 365218
rect 92114 331538 92146 331774
rect 92382 331538 92466 331774
rect 92702 331538 92734 331774
rect 92114 331454 92734 331538
rect 92114 331218 92146 331454
rect 92382 331218 92466 331454
rect 92702 331218 92734 331454
rect 92114 297774 92734 331218
rect 92114 297538 92146 297774
rect 92382 297538 92466 297774
rect 92702 297538 92734 297774
rect 92114 297454 92734 297538
rect 92114 297218 92146 297454
rect 92382 297218 92466 297454
rect 92702 297218 92734 297454
rect 92114 263774 92734 297218
rect 92114 263538 92146 263774
rect 92382 263538 92466 263774
rect 92702 263538 92734 263774
rect 92114 263454 92734 263538
rect 92114 263218 92146 263454
rect 92382 263218 92466 263454
rect 92702 263218 92734 263454
rect 92114 229774 92734 263218
rect 92114 229538 92146 229774
rect 92382 229538 92466 229774
rect 92702 229538 92734 229774
rect 92114 229454 92734 229538
rect 92114 229218 92146 229454
rect 92382 229218 92466 229454
rect 92702 229218 92734 229454
rect 92114 225660 92734 229218
rect 95834 711558 96454 711590
rect 95834 711322 95866 711558
rect 96102 711322 96186 711558
rect 96422 711322 96454 711558
rect 95834 711238 96454 711322
rect 95834 711002 95866 711238
rect 96102 711002 96186 711238
rect 96422 711002 96454 711238
rect 95834 675494 96454 711002
rect 95834 675258 95866 675494
rect 96102 675258 96186 675494
rect 96422 675258 96454 675494
rect 95834 675174 96454 675258
rect 95834 674938 95866 675174
rect 96102 674938 96186 675174
rect 96422 674938 96454 675174
rect 95834 641494 96454 674938
rect 95834 641258 95866 641494
rect 96102 641258 96186 641494
rect 96422 641258 96454 641494
rect 95834 641174 96454 641258
rect 95834 640938 95866 641174
rect 96102 640938 96186 641174
rect 96422 640938 96454 641174
rect 95834 607494 96454 640938
rect 95834 607258 95866 607494
rect 96102 607258 96186 607494
rect 96422 607258 96454 607494
rect 95834 607174 96454 607258
rect 95834 606938 95866 607174
rect 96102 606938 96186 607174
rect 96422 606938 96454 607174
rect 95834 573494 96454 606938
rect 95834 573258 95866 573494
rect 96102 573258 96186 573494
rect 96422 573258 96454 573494
rect 95834 573174 96454 573258
rect 95834 572938 95866 573174
rect 96102 572938 96186 573174
rect 96422 572938 96454 573174
rect 95834 539494 96454 572938
rect 95834 539258 95866 539494
rect 96102 539258 96186 539494
rect 96422 539258 96454 539494
rect 95834 539174 96454 539258
rect 95834 538938 95866 539174
rect 96102 538938 96186 539174
rect 96422 538938 96454 539174
rect 95834 505494 96454 538938
rect 95834 505258 95866 505494
rect 96102 505258 96186 505494
rect 96422 505258 96454 505494
rect 95834 505174 96454 505258
rect 95834 504938 95866 505174
rect 96102 504938 96186 505174
rect 96422 504938 96454 505174
rect 95834 471494 96454 504938
rect 95834 471258 95866 471494
rect 96102 471258 96186 471494
rect 96422 471258 96454 471494
rect 95834 471174 96454 471258
rect 95834 470938 95866 471174
rect 96102 470938 96186 471174
rect 96422 470938 96454 471174
rect 95834 437494 96454 470938
rect 95834 437258 95866 437494
rect 96102 437258 96186 437494
rect 96422 437258 96454 437494
rect 95834 437174 96454 437258
rect 95834 436938 95866 437174
rect 96102 436938 96186 437174
rect 96422 436938 96454 437174
rect 95834 403494 96454 436938
rect 95834 403258 95866 403494
rect 96102 403258 96186 403494
rect 96422 403258 96454 403494
rect 95834 403174 96454 403258
rect 95834 402938 95866 403174
rect 96102 402938 96186 403174
rect 96422 402938 96454 403174
rect 95834 369494 96454 402938
rect 95834 369258 95866 369494
rect 96102 369258 96186 369494
rect 96422 369258 96454 369494
rect 95834 369174 96454 369258
rect 95834 368938 95866 369174
rect 96102 368938 96186 369174
rect 96422 368938 96454 369174
rect 95834 335494 96454 368938
rect 95834 335258 95866 335494
rect 96102 335258 96186 335494
rect 96422 335258 96454 335494
rect 95834 335174 96454 335258
rect 95834 334938 95866 335174
rect 96102 334938 96186 335174
rect 96422 334938 96454 335174
rect 95834 301494 96454 334938
rect 95834 301258 95866 301494
rect 96102 301258 96186 301494
rect 96422 301258 96454 301494
rect 95834 301174 96454 301258
rect 95834 300938 95866 301174
rect 96102 300938 96186 301174
rect 96422 300938 96454 301174
rect 95834 267494 96454 300938
rect 95834 267258 95866 267494
rect 96102 267258 96186 267494
rect 96422 267258 96454 267494
rect 95834 267174 96454 267258
rect 95834 266938 95866 267174
rect 96102 266938 96186 267174
rect 96422 266938 96454 267174
rect 95834 233494 96454 266938
rect 95834 233258 95866 233494
rect 96102 233258 96186 233494
rect 96422 233258 96454 233494
rect 95834 233174 96454 233258
rect 95834 232938 95866 233174
rect 96102 232938 96186 233174
rect 96422 232938 96454 233174
rect 95834 225660 96454 232938
rect 103794 704838 104414 711590
rect 103794 704602 103826 704838
rect 104062 704602 104146 704838
rect 104382 704602 104414 704838
rect 103794 704518 104414 704602
rect 103794 704282 103826 704518
rect 104062 704282 104146 704518
rect 104382 704282 104414 704518
rect 103794 683454 104414 704282
rect 103794 683218 103826 683454
rect 104062 683218 104146 683454
rect 104382 683218 104414 683454
rect 103794 683134 104414 683218
rect 103794 682898 103826 683134
rect 104062 682898 104146 683134
rect 104382 682898 104414 683134
rect 103794 649454 104414 682898
rect 103794 649218 103826 649454
rect 104062 649218 104146 649454
rect 104382 649218 104414 649454
rect 103794 649134 104414 649218
rect 103794 648898 103826 649134
rect 104062 648898 104146 649134
rect 104382 648898 104414 649134
rect 103794 615454 104414 648898
rect 103794 615218 103826 615454
rect 104062 615218 104146 615454
rect 104382 615218 104414 615454
rect 103794 615134 104414 615218
rect 103794 614898 103826 615134
rect 104062 614898 104146 615134
rect 104382 614898 104414 615134
rect 103794 581454 104414 614898
rect 103794 581218 103826 581454
rect 104062 581218 104146 581454
rect 104382 581218 104414 581454
rect 103794 581134 104414 581218
rect 103794 580898 103826 581134
rect 104062 580898 104146 581134
rect 104382 580898 104414 581134
rect 103794 547454 104414 580898
rect 103794 547218 103826 547454
rect 104062 547218 104146 547454
rect 104382 547218 104414 547454
rect 103794 547134 104414 547218
rect 103794 546898 103826 547134
rect 104062 546898 104146 547134
rect 104382 546898 104414 547134
rect 103794 513454 104414 546898
rect 103794 513218 103826 513454
rect 104062 513218 104146 513454
rect 104382 513218 104414 513454
rect 103794 513134 104414 513218
rect 103794 512898 103826 513134
rect 104062 512898 104146 513134
rect 104382 512898 104414 513134
rect 103794 479454 104414 512898
rect 103794 479218 103826 479454
rect 104062 479218 104146 479454
rect 104382 479218 104414 479454
rect 103794 479134 104414 479218
rect 103794 478898 103826 479134
rect 104062 478898 104146 479134
rect 104382 478898 104414 479134
rect 103794 445454 104414 478898
rect 103794 445218 103826 445454
rect 104062 445218 104146 445454
rect 104382 445218 104414 445454
rect 103794 445134 104414 445218
rect 103794 444898 103826 445134
rect 104062 444898 104146 445134
rect 104382 444898 104414 445134
rect 103794 411454 104414 444898
rect 103794 411218 103826 411454
rect 104062 411218 104146 411454
rect 104382 411218 104414 411454
rect 103794 411134 104414 411218
rect 103794 410898 103826 411134
rect 104062 410898 104146 411134
rect 104382 410898 104414 411134
rect 103794 377454 104414 410898
rect 103794 377218 103826 377454
rect 104062 377218 104146 377454
rect 104382 377218 104414 377454
rect 103794 377134 104414 377218
rect 103794 376898 103826 377134
rect 104062 376898 104146 377134
rect 104382 376898 104414 377134
rect 103794 343454 104414 376898
rect 103794 343218 103826 343454
rect 104062 343218 104146 343454
rect 104382 343218 104414 343454
rect 103794 343134 104414 343218
rect 103794 342898 103826 343134
rect 104062 342898 104146 343134
rect 104382 342898 104414 343134
rect 103794 309454 104414 342898
rect 103794 309218 103826 309454
rect 104062 309218 104146 309454
rect 104382 309218 104414 309454
rect 103794 309134 104414 309218
rect 103794 308898 103826 309134
rect 104062 308898 104146 309134
rect 104382 308898 104414 309134
rect 103794 275454 104414 308898
rect 103794 275218 103826 275454
rect 104062 275218 104146 275454
rect 104382 275218 104414 275454
rect 103794 275134 104414 275218
rect 103794 274898 103826 275134
rect 104062 274898 104146 275134
rect 104382 274898 104414 275134
rect 103794 241454 104414 274898
rect 103794 241218 103826 241454
rect 104062 241218 104146 241454
rect 104382 241218 104414 241454
rect 103794 241134 104414 241218
rect 103794 240898 103826 241134
rect 104062 240898 104146 241134
rect 104382 240898 104414 241134
rect 103794 225660 104414 240898
rect 107514 705798 108134 711590
rect 107514 705562 107546 705798
rect 107782 705562 107866 705798
rect 108102 705562 108134 705798
rect 107514 705478 108134 705562
rect 107514 705242 107546 705478
rect 107782 705242 107866 705478
rect 108102 705242 108134 705478
rect 107514 687174 108134 705242
rect 107514 686938 107546 687174
rect 107782 686938 107866 687174
rect 108102 686938 108134 687174
rect 107514 686854 108134 686938
rect 107514 686618 107546 686854
rect 107782 686618 107866 686854
rect 108102 686618 108134 686854
rect 107514 653174 108134 686618
rect 107514 652938 107546 653174
rect 107782 652938 107866 653174
rect 108102 652938 108134 653174
rect 107514 652854 108134 652938
rect 107514 652618 107546 652854
rect 107782 652618 107866 652854
rect 108102 652618 108134 652854
rect 107514 619174 108134 652618
rect 107514 618938 107546 619174
rect 107782 618938 107866 619174
rect 108102 618938 108134 619174
rect 107514 618854 108134 618938
rect 107514 618618 107546 618854
rect 107782 618618 107866 618854
rect 108102 618618 108134 618854
rect 107514 585174 108134 618618
rect 107514 584938 107546 585174
rect 107782 584938 107866 585174
rect 108102 584938 108134 585174
rect 107514 584854 108134 584938
rect 107514 584618 107546 584854
rect 107782 584618 107866 584854
rect 108102 584618 108134 584854
rect 107514 551174 108134 584618
rect 107514 550938 107546 551174
rect 107782 550938 107866 551174
rect 108102 550938 108134 551174
rect 107514 550854 108134 550938
rect 107514 550618 107546 550854
rect 107782 550618 107866 550854
rect 108102 550618 108134 550854
rect 107514 517174 108134 550618
rect 107514 516938 107546 517174
rect 107782 516938 107866 517174
rect 108102 516938 108134 517174
rect 107514 516854 108134 516938
rect 107514 516618 107546 516854
rect 107782 516618 107866 516854
rect 108102 516618 108134 516854
rect 107514 483174 108134 516618
rect 107514 482938 107546 483174
rect 107782 482938 107866 483174
rect 108102 482938 108134 483174
rect 107514 482854 108134 482938
rect 107514 482618 107546 482854
rect 107782 482618 107866 482854
rect 108102 482618 108134 482854
rect 107514 449174 108134 482618
rect 107514 448938 107546 449174
rect 107782 448938 107866 449174
rect 108102 448938 108134 449174
rect 107514 448854 108134 448938
rect 107514 448618 107546 448854
rect 107782 448618 107866 448854
rect 108102 448618 108134 448854
rect 107514 415174 108134 448618
rect 107514 414938 107546 415174
rect 107782 414938 107866 415174
rect 108102 414938 108134 415174
rect 107514 414854 108134 414938
rect 107514 414618 107546 414854
rect 107782 414618 107866 414854
rect 108102 414618 108134 414854
rect 107514 381174 108134 414618
rect 107514 380938 107546 381174
rect 107782 380938 107866 381174
rect 108102 380938 108134 381174
rect 107514 380854 108134 380938
rect 107514 380618 107546 380854
rect 107782 380618 107866 380854
rect 108102 380618 108134 380854
rect 107514 347174 108134 380618
rect 107514 346938 107546 347174
rect 107782 346938 107866 347174
rect 108102 346938 108134 347174
rect 107514 346854 108134 346938
rect 107514 346618 107546 346854
rect 107782 346618 107866 346854
rect 108102 346618 108134 346854
rect 107514 313174 108134 346618
rect 107514 312938 107546 313174
rect 107782 312938 107866 313174
rect 108102 312938 108134 313174
rect 107514 312854 108134 312938
rect 107514 312618 107546 312854
rect 107782 312618 107866 312854
rect 108102 312618 108134 312854
rect 107514 279174 108134 312618
rect 107514 278938 107546 279174
rect 107782 278938 107866 279174
rect 108102 278938 108134 279174
rect 107514 278854 108134 278938
rect 107514 278618 107546 278854
rect 107782 278618 107866 278854
rect 108102 278618 108134 278854
rect 107514 245174 108134 278618
rect 107514 244938 107546 245174
rect 107782 244938 107866 245174
rect 108102 244938 108134 245174
rect 107514 244854 108134 244938
rect 107514 244618 107546 244854
rect 107782 244618 107866 244854
rect 108102 244618 108134 244854
rect 107514 225660 108134 244618
rect 111234 706758 111854 711590
rect 111234 706522 111266 706758
rect 111502 706522 111586 706758
rect 111822 706522 111854 706758
rect 111234 706438 111854 706522
rect 111234 706202 111266 706438
rect 111502 706202 111586 706438
rect 111822 706202 111854 706438
rect 111234 690894 111854 706202
rect 111234 690658 111266 690894
rect 111502 690658 111586 690894
rect 111822 690658 111854 690894
rect 111234 690574 111854 690658
rect 111234 690338 111266 690574
rect 111502 690338 111586 690574
rect 111822 690338 111854 690574
rect 111234 656894 111854 690338
rect 111234 656658 111266 656894
rect 111502 656658 111586 656894
rect 111822 656658 111854 656894
rect 111234 656574 111854 656658
rect 111234 656338 111266 656574
rect 111502 656338 111586 656574
rect 111822 656338 111854 656574
rect 111234 622894 111854 656338
rect 111234 622658 111266 622894
rect 111502 622658 111586 622894
rect 111822 622658 111854 622894
rect 111234 622574 111854 622658
rect 111234 622338 111266 622574
rect 111502 622338 111586 622574
rect 111822 622338 111854 622574
rect 111234 588894 111854 622338
rect 111234 588658 111266 588894
rect 111502 588658 111586 588894
rect 111822 588658 111854 588894
rect 111234 588574 111854 588658
rect 111234 588338 111266 588574
rect 111502 588338 111586 588574
rect 111822 588338 111854 588574
rect 111234 554894 111854 588338
rect 111234 554658 111266 554894
rect 111502 554658 111586 554894
rect 111822 554658 111854 554894
rect 111234 554574 111854 554658
rect 111234 554338 111266 554574
rect 111502 554338 111586 554574
rect 111822 554338 111854 554574
rect 111234 520894 111854 554338
rect 111234 520658 111266 520894
rect 111502 520658 111586 520894
rect 111822 520658 111854 520894
rect 111234 520574 111854 520658
rect 111234 520338 111266 520574
rect 111502 520338 111586 520574
rect 111822 520338 111854 520574
rect 111234 486894 111854 520338
rect 111234 486658 111266 486894
rect 111502 486658 111586 486894
rect 111822 486658 111854 486894
rect 111234 486574 111854 486658
rect 111234 486338 111266 486574
rect 111502 486338 111586 486574
rect 111822 486338 111854 486574
rect 111234 452894 111854 486338
rect 111234 452658 111266 452894
rect 111502 452658 111586 452894
rect 111822 452658 111854 452894
rect 111234 452574 111854 452658
rect 111234 452338 111266 452574
rect 111502 452338 111586 452574
rect 111822 452338 111854 452574
rect 111234 418894 111854 452338
rect 111234 418658 111266 418894
rect 111502 418658 111586 418894
rect 111822 418658 111854 418894
rect 111234 418574 111854 418658
rect 111234 418338 111266 418574
rect 111502 418338 111586 418574
rect 111822 418338 111854 418574
rect 111234 384894 111854 418338
rect 111234 384658 111266 384894
rect 111502 384658 111586 384894
rect 111822 384658 111854 384894
rect 111234 384574 111854 384658
rect 111234 384338 111266 384574
rect 111502 384338 111586 384574
rect 111822 384338 111854 384574
rect 111234 350894 111854 384338
rect 111234 350658 111266 350894
rect 111502 350658 111586 350894
rect 111822 350658 111854 350894
rect 111234 350574 111854 350658
rect 111234 350338 111266 350574
rect 111502 350338 111586 350574
rect 111822 350338 111854 350574
rect 111234 316894 111854 350338
rect 111234 316658 111266 316894
rect 111502 316658 111586 316894
rect 111822 316658 111854 316894
rect 111234 316574 111854 316658
rect 111234 316338 111266 316574
rect 111502 316338 111586 316574
rect 111822 316338 111854 316574
rect 111234 282894 111854 316338
rect 111234 282658 111266 282894
rect 111502 282658 111586 282894
rect 111822 282658 111854 282894
rect 111234 282574 111854 282658
rect 111234 282338 111266 282574
rect 111502 282338 111586 282574
rect 111822 282338 111854 282574
rect 111234 248894 111854 282338
rect 111234 248658 111266 248894
rect 111502 248658 111586 248894
rect 111822 248658 111854 248894
rect 111234 248574 111854 248658
rect 111234 248338 111266 248574
rect 111502 248338 111586 248574
rect 111822 248338 111854 248574
rect 111234 225660 111854 248338
rect 114954 707718 115574 711590
rect 114954 707482 114986 707718
rect 115222 707482 115306 707718
rect 115542 707482 115574 707718
rect 114954 707398 115574 707482
rect 114954 707162 114986 707398
rect 115222 707162 115306 707398
rect 115542 707162 115574 707398
rect 114954 694614 115574 707162
rect 114954 694378 114986 694614
rect 115222 694378 115306 694614
rect 115542 694378 115574 694614
rect 114954 694294 115574 694378
rect 114954 694058 114986 694294
rect 115222 694058 115306 694294
rect 115542 694058 115574 694294
rect 114954 660614 115574 694058
rect 114954 660378 114986 660614
rect 115222 660378 115306 660614
rect 115542 660378 115574 660614
rect 114954 660294 115574 660378
rect 114954 660058 114986 660294
rect 115222 660058 115306 660294
rect 115542 660058 115574 660294
rect 114954 626614 115574 660058
rect 114954 626378 114986 626614
rect 115222 626378 115306 626614
rect 115542 626378 115574 626614
rect 114954 626294 115574 626378
rect 114954 626058 114986 626294
rect 115222 626058 115306 626294
rect 115542 626058 115574 626294
rect 114954 592614 115574 626058
rect 114954 592378 114986 592614
rect 115222 592378 115306 592614
rect 115542 592378 115574 592614
rect 114954 592294 115574 592378
rect 114954 592058 114986 592294
rect 115222 592058 115306 592294
rect 115542 592058 115574 592294
rect 114954 558614 115574 592058
rect 114954 558378 114986 558614
rect 115222 558378 115306 558614
rect 115542 558378 115574 558614
rect 114954 558294 115574 558378
rect 114954 558058 114986 558294
rect 115222 558058 115306 558294
rect 115542 558058 115574 558294
rect 114954 524614 115574 558058
rect 114954 524378 114986 524614
rect 115222 524378 115306 524614
rect 115542 524378 115574 524614
rect 114954 524294 115574 524378
rect 114954 524058 114986 524294
rect 115222 524058 115306 524294
rect 115542 524058 115574 524294
rect 114954 490614 115574 524058
rect 114954 490378 114986 490614
rect 115222 490378 115306 490614
rect 115542 490378 115574 490614
rect 114954 490294 115574 490378
rect 114954 490058 114986 490294
rect 115222 490058 115306 490294
rect 115542 490058 115574 490294
rect 114954 456614 115574 490058
rect 114954 456378 114986 456614
rect 115222 456378 115306 456614
rect 115542 456378 115574 456614
rect 114954 456294 115574 456378
rect 114954 456058 114986 456294
rect 115222 456058 115306 456294
rect 115542 456058 115574 456294
rect 114954 422614 115574 456058
rect 114954 422378 114986 422614
rect 115222 422378 115306 422614
rect 115542 422378 115574 422614
rect 114954 422294 115574 422378
rect 114954 422058 114986 422294
rect 115222 422058 115306 422294
rect 115542 422058 115574 422294
rect 114954 388614 115574 422058
rect 114954 388378 114986 388614
rect 115222 388378 115306 388614
rect 115542 388378 115574 388614
rect 114954 388294 115574 388378
rect 114954 388058 114986 388294
rect 115222 388058 115306 388294
rect 115542 388058 115574 388294
rect 114954 354614 115574 388058
rect 114954 354378 114986 354614
rect 115222 354378 115306 354614
rect 115542 354378 115574 354614
rect 114954 354294 115574 354378
rect 114954 354058 114986 354294
rect 115222 354058 115306 354294
rect 115542 354058 115574 354294
rect 114954 320614 115574 354058
rect 114954 320378 114986 320614
rect 115222 320378 115306 320614
rect 115542 320378 115574 320614
rect 114954 320294 115574 320378
rect 114954 320058 114986 320294
rect 115222 320058 115306 320294
rect 115542 320058 115574 320294
rect 114954 286614 115574 320058
rect 114954 286378 114986 286614
rect 115222 286378 115306 286614
rect 115542 286378 115574 286614
rect 114954 286294 115574 286378
rect 114954 286058 114986 286294
rect 115222 286058 115306 286294
rect 115542 286058 115574 286294
rect 114954 252614 115574 286058
rect 114954 252378 114986 252614
rect 115222 252378 115306 252614
rect 115542 252378 115574 252614
rect 114954 252294 115574 252378
rect 114954 252058 114986 252294
rect 115222 252058 115306 252294
rect 115542 252058 115574 252294
rect 114954 225660 115574 252058
rect 118674 708678 119294 711590
rect 118674 708442 118706 708678
rect 118942 708442 119026 708678
rect 119262 708442 119294 708678
rect 118674 708358 119294 708442
rect 118674 708122 118706 708358
rect 118942 708122 119026 708358
rect 119262 708122 119294 708358
rect 118674 698334 119294 708122
rect 118674 698098 118706 698334
rect 118942 698098 119026 698334
rect 119262 698098 119294 698334
rect 118674 698014 119294 698098
rect 118674 697778 118706 698014
rect 118942 697778 119026 698014
rect 119262 697778 119294 698014
rect 118674 664334 119294 697778
rect 118674 664098 118706 664334
rect 118942 664098 119026 664334
rect 119262 664098 119294 664334
rect 118674 664014 119294 664098
rect 118674 663778 118706 664014
rect 118942 663778 119026 664014
rect 119262 663778 119294 664014
rect 118674 630334 119294 663778
rect 118674 630098 118706 630334
rect 118942 630098 119026 630334
rect 119262 630098 119294 630334
rect 118674 630014 119294 630098
rect 118674 629778 118706 630014
rect 118942 629778 119026 630014
rect 119262 629778 119294 630014
rect 118674 596334 119294 629778
rect 118674 596098 118706 596334
rect 118942 596098 119026 596334
rect 119262 596098 119294 596334
rect 118674 596014 119294 596098
rect 118674 595778 118706 596014
rect 118942 595778 119026 596014
rect 119262 595778 119294 596014
rect 118674 562334 119294 595778
rect 118674 562098 118706 562334
rect 118942 562098 119026 562334
rect 119262 562098 119294 562334
rect 118674 562014 119294 562098
rect 118674 561778 118706 562014
rect 118942 561778 119026 562014
rect 119262 561778 119294 562014
rect 118674 528334 119294 561778
rect 118674 528098 118706 528334
rect 118942 528098 119026 528334
rect 119262 528098 119294 528334
rect 118674 528014 119294 528098
rect 118674 527778 118706 528014
rect 118942 527778 119026 528014
rect 119262 527778 119294 528014
rect 118674 494334 119294 527778
rect 118674 494098 118706 494334
rect 118942 494098 119026 494334
rect 119262 494098 119294 494334
rect 118674 494014 119294 494098
rect 118674 493778 118706 494014
rect 118942 493778 119026 494014
rect 119262 493778 119294 494014
rect 118674 460334 119294 493778
rect 118674 460098 118706 460334
rect 118942 460098 119026 460334
rect 119262 460098 119294 460334
rect 118674 460014 119294 460098
rect 118674 459778 118706 460014
rect 118942 459778 119026 460014
rect 119262 459778 119294 460014
rect 118674 426334 119294 459778
rect 118674 426098 118706 426334
rect 118942 426098 119026 426334
rect 119262 426098 119294 426334
rect 118674 426014 119294 426098
rect 118674 425778 118706 426014
rect 118942 425778 119026 426014
rect 119262 425778 119294 426014
rect 118674 392334 119294 425778
rect 118674 392098 118706 392334
rect 118942 392098 119026 392334
rect 119262 392098 119294 392334
rect 118674 392014 119294 392098
rect 118674 391778 118706 392014
rect 118942 391778 119026 392014
rect 119262 391778 119294 392014
rect 118674 358334 119294 391778
rect 118674 358098 118706 358334
rect 118942 358098 119026 358334
rect 119262 358098 119294 358334
rect 118674 358014 119294 358098
rect 118674 357778 118706 358014
rect 118942 357778 119026 358014
rect 119262 357778 119294 358014
rect 118674 324334 119294 357778
rect 118674 324098 118706 324334
rect 118942 324098 119026 324334
rect 119262 324098 119294 324334
rect 118674 324014 119294 324098
rect 118674 323778 118706 324014
rect 118942 323778 119026 324014
rect 119262 323778 119294 324014
rect 118674 290334 119294 323778
rect 118674 290098 118706 290334
rect 118942 290098 119026 290334
rect 119262 290098 119294 290334
rect 118674 290014 119294 290098
rect 118674 289778 118706 290014
rect 118942 289778 119026 290014
rect 119262 289778 119294 290014
rect 118674 256334 119294 289778
rect 118674 256098 118706 256334
rect 118942 256098 119026 256334
rect 119262 256098 119294 256334
rect 118674 256014 119294 256098
rect 118674 255778 118706 256014
rect 118942 255778 119026 256014
rect 119262 255778 119294 256014
rect 118674 225660 119294 255778
rect 122394 709638 123014 711590
rect 122394 709402 122426 709638
rect 122662 709402 122746 709638
rect 122982 709402 123014 709638
rect 122394 709318 123014 709402
rect 122394 709082 122426 709318
rect 122662 709082 122746 709318
rect 122982 709082 123014 709318
rect 122394 668054 123014 709082
rect 122394 667818 122426 668054
rect 122662 667818 122746 668054
rect 122982 667818 123014 668054
rect 122394 667734 123014 667818
rect 122394 667498 122426 667734
rect 122662 667498 122746 667734
rect 122982 667498 123014 667734
rect 122394 634054 123014 667498
rect 122394 633818 122426 634054
rect 122662 633818 122746 634054
rect 122982 633818 123014 634054
rect 122394 633734 123014 633818
rect 122394 633498 122426 633734
rect 122662 633498 122746 633734
rect 122982 633498 123014 633734
rect 122394 600054 123014 633498
rect 122394 599818 122426 600054
rect 122662 599818 122746 600054
rect 122982 599818 123014 600054
rect 122394 599734 123014 599818
rect 122394 599498 122426 599734
rect 122662 599498 122746 599734
rect 122982 599498 123014 599734
rect 122394 566054 123014 599498
rect 122394 565818 122426 566054
rect 122662 565818 122746 566054
rect 122982 565818 123014 566054
rect 122394 565734 123014 565818
rect 122394 565498 122426 565734
rect 122662 565498 122746 565734
rect 122982 565498 123014 565734
rect 122394 532054 123014 565498
rect 122394 531818 122426 532054
rect 122662 531818 122746 532054
rect 122982 531818 123014 532054
rect 122394 531734 123014 531818
rect 122394 531498 122426 531734
rect 122662 531498 122746 531734
rect 122982 531498 123014 531734
rect 122394 498054 123014 531498
rect 122394 497818 122426 498054
rect 122662 497818 122746 498054
rect 122982 497818 123014 498054
rect 122394 497734 123014 497818
rect 122394 497498 122426 497734
rect 122662 497498 122746 497734
rect 122982 497498 123014 497734
rect 122394 464054 123014 497498
rect 122394 463818 122426 464054
rect 122662 463818 122746 464054
rect 122982 463818 123014 464054
rect 122394 463734 123014 463818
rect 122394 463498 122426 463734
rect 122662 463498 122746 463734
rect 122982 463498 123014 463734
rect 122394 430054 123014 463498
rect 122394 429818 122426 430054
rect 122662 429818 122746 430054
rect 122982 429818 123014 430054
rect 122394 429734 123014 429818
rect 122394 429498 122426 429734
rect 122662 429498 122746 429734
rect 122982 429498 123014 429734
rect 122394 396054 123014 429498
rect 122394 395818 122426 396054
rect 122662 395818 122746 396054
rect 122982 395818 123014 396054
rect 122394 395734 123014 395818
rect 122394 395498 122426 395734
rect 122662 395498 122746 395734
rect 122982 395498 123014 395734
rect 122394 362054 123014 395498
rect 122394 361818 122426 362054
rect 122662 361818 122746 362054
rect 122982 361818 123014 362054
rect 122394 361734 123014 361818
rect 122394 361498 122426 361734
rect 122662 361498 122746 361734
rect 122982 361498 123014 361734
rect 122394 328054 123014 361498
rect 122394 327818 122426 328054
rect 122662 327818 122746 328054
rect 122982 327818 123014 328054
rect 122394 327734 123014 327818
rect 122394 327498 122426 327734
rect 122662 327498 122746 327734
rect 122982 327498 123014 327734
rect 122394 294054 123014 327498
rect 122394 293818 122426 294054
rect 122662 293818 122746 294054
rect 122982 293818 123014 294054
rect 122394 293734 123014 293818
rect 122394 293498 122426 293734
rect 122662 293498 122746 293734
rect 122982 293498 123014 293734
rect 122394 260054 123014 293498
rect 122394 259818 122426 260054
rect 122662 259818 122746 260054
rect 122982 259818 123014 260054
rect 122394 259734 123014 259818
rect 122394 259498 122426 259734
rect 122662 259498 122746 259734
rect 122982 259498 123014 259734
rect 122394 225991 123014 259498
rect 122394 225755 122426 225991
rect 122662 225755 122746 225991
rect 122982 225755 123014 225991
rect 122394 225660 123014 225755
rect 126114 710598 126734 711590
rect 126114 710362 126146 710598
rect 126382 710362 126466 710598
rect 126702 710362 126734 710598
rect 126114 710278 126734 710362
rect 126114 710042 126146 710278
rect 126382 710042 126466 710278
rect 126702 710042 126734 710278
rect 126114 671774 126734 710042
rect 126114 671538 126146 671774
rect 126382 671538 126466 671774
rect 126702 671538 126734 671774
rect 126114 671454 126734 671538
rect 126114 671218 126146 671454
rect 126382 671218 126466 671454
rect 126702 671218 126734 671454
rect 126114 637774 126734 671218
rect 126114 637538 126146 637774
rect 126382 637538 126466 637774
rect 126702 637538 126734 637774
rect 126114 637454 126734 637538
rect 126114 637218 126146 637454
rect 126382 637218 126466 637454
rect 126702 637218 126734 637454
rect 126114 603774 126734 637218
rect 126114 603538 126146 603774
rect 126382 603538 126466 603774
rect 126702 603538 126734 603774
rect 126114 603454 126734 603538
rect 126114 603218 126146 603454
rect 126382 603218 126466 603454
rect 126702 603218 126734 603454
rect 126114 569774 126734 603218
rect 126114 569538 126146 569774
rect 126382 569538 126466 569774
rect 126702 569538 126734 569774
rect 126114 569454 126734 569538
rect 126114 569218 126146 569454
rect 126382 569218 126466 569454
rect 126702 569218 126734 569454
rect 126114 535774 126734 569218
rect 126114 535538 126146 535774
rect 126382 535538 126466 535774
rect 126702 535538 126734 535774
rect 126114 535454 126734 535538
rect 126114 535218 126146 535454
rect 126382 535218 126466 535454
rect 126702 535218 126734 535454
rect 126114 501774 126734 535218
rect 126114 501538 126146 501774
rect 126382 501538 126466 501774
rect 126702 501538 126734 501774
rect 126114 501454 126734 501538
rect 126114 501218 126146 501454
rect 126382 501218 126466 501454
rect 126702 501218 126734 501454
rect 126114 467774 126734 501218
rect 126114 467538 126146 467774
rect 126382 467538 126466 467774
rect 126702 467538 126734 467774
rect 126114 467454 126734 467538
rect 126114 467218 126146 467454
rect 126382 467218 126466 467454
rect 126702 467218 126734 467454
rect 126114 433774 126734 467218
rect 126114 433538 126146 433774
rect 126382 433538 126466 433774
rect 126702 433538 126734 433774
rect 126114 433454 126734 433538
rect 126114 433218 126146 433454
rect 126382 433218 126466 433454
rect 126702 433218 126734 433454
rect 126114 399774 126734 433218
rect 126114 399538 126146 399774
rect 126382 399538 126466 399774
rect 126702 399538 126734 399774
rect 126114 399454 126734 399538
rect 126114 399218 126146 399454
rect 126382 399218 126466 399454
rect 126702 399218 126734 399454
rect 126114 365774 126734 399218
rect 126114 365538 126146 365774
rect 126382 365538 126466 365774
rect 126702 365538 126734 365774
rect 126114 365454 126734 365538
rect 126114 365218 126146 365454
rect 126382 365218 126466 365454
rect 126702 365218 126734 365454
rect 126114 331774 126734 365218
rect 126114 331538 126146 331774
rect 126382 331538 126466 331774
rect 126702 331538 126734 331774
rect 126114 331454 126734 331538
rect 126114 331218 126146 331454
rect 126382 331218 126466 331454
rect 126702 331218 126734 331454
rect 126114 297774 126734 331218
rect 126114 297538 126146 297774
rect 126382 297538 126466 297774
rect 126702 297538 126734 297774
rect 126114 297454 126734 297538
rect 126114 297218 126146 297454
rect 126382 297218 126466 297454
rect 126702 297218 126734 297454
rect 126114 263774 126734 297218
rect 126114 263538 126146 263774
rect 126382 263538 126466 263774
rect 126702 263538 126734 263774
rect 126114 263454 126734 263538
rect 126114 263218 126146 263454
rect 126382 263218 126466 263454
rect 126702 263218 126734 263454
rect 126114 229774 126734 263218
rect 126114 229538 126146 229774
rect 126382 229538 126466 229774
rect 126702 229538 126734 229774
rect 126114 229454 126734 229538
rect 126114 229218 126146 229454
rect 126382 229218 126466 229454
rect 126702 229218 126734 229454
rect 126114 225660 126734 229218
rect 129834 711558 130454 711590
rect 129834 711322 129866 711558
rect 130102 711322 130186 711558
rect 130422 711322 130454 711558
rect 129834 711238 130454 711322
rect 129834 711002 129866 711238
rect 130102 711002 130186 711238
rect 130422 711002 130454 711238
rect 129834 675494 130454 711002
rect 129834 675258 129866 675494
rect 130102 675258 130186 675494
rect 130422 675258 130454 675494
rect 129834 675174 130454 675258
rect 129834 674938 129866 675174
rect 130102 674938 130186 675174
rect 130422 674938 130454 675174
rect 129834 641494 130454 674938
rect 129834 641258 129866 641494
rect 130102 641258 130186 641494
rect 130422 641258 130454 641494
rect 129834 641174 130454 641258
rect 129834 640938 129866 641174
rect 130102 640938 130186 641174
rect 130422 640938 130454 641174
rect 129834 607494 130454 640938
rect 129834 607258 129866 607494
rect 130102 607258 130186 607494
rect 130422 607258 130454 607494
rect 129834 607174 130454 607258
rect 129834 606938 129866 607174
rect 130102 606938 130186 607174
rect 130422 606938 130454 607174
rect 129834 573494 130454 606938
rect 129834 573258 129866 573494
rect 130102 573258 130186 573494
rect 130422 573258 130454 573494
rect 129834 573174 130454 573258
rect 129834 572938 129866 573174
rect 130102 572938 130186 573174
rect 130422 572938 130454 573174
rect 129834 539494 130454 572938
rect 129834 539258 129866 539494
rect 130102 539258 130186 539494
rect 130422 539258 130454 539494
rect 129834 539174 130454 539258
rect 129834 538938 129866 539174
rect 130102 538938 130186 539174
rect 130422 538938 130454 539174
rect 129834 505494 130454 538938
rect 129834 505258 129866 505494
rect 130102 505258 130186 505494
rect 130422 505258 130454 505494
rect 129834 505174 130454 505258
rect 129834 504938 129866 505174
rect 130102 504938 130186 505174
rect 130422 504938 130454 505174
rect 129834 471494 130454 504938
rect 129834 471258 129866 471494
rect 130102 471258 130186 471494
rect 130422 471258 130454 471494
rect 129834 471174 130454 471258
rect 129834 470938 129866 471174
rect 130102 470938 130186 471174
rect 130422 470938 130454 471174
rect 129834 437494 130454 470938
rect 129834 437258 129866 437494
rect 130102 437258 130186 437494
rect 130422 437258 130454 437494
rect 129834 437174 130454 437258
rect 129834 436938 129866 437174
rect 130102 436938 130186 437174
rect 130422 436938 130454 437174
rect 129834 403494 130454 436938
rect 129834 403258 129866 403494
rect 130102 403258 130186 403494
rect 130422 403258 130454 403494
rect 129834 403174 130454 403258
rect 129834 402938 129866 403174
rect 130102 402938 130186 403174
rect 130422 402938 130454 403174
rect 129834 369494 130454 402938
rect 129834 369258 129866 369494
rect 130102 369258 130186 369494
rect 130422 369258 130454 369494
rect 129834 369174 130454 369258
rect 129834 368938 129866 369174
rect 130102 368938 130186 369174
rect 130422 368938 130454 369174
rect 129834 335494 130454 368938
rect 129834 335258 129866 335494
rect 130102 335258 130186 335494
rect 130422 335258 130454 335494
rect 129834 335174 130454 335258
rect 129834 334938 129866 335174
rect 130102 334938 130186 335174
rect 130422 334938 130454 335174
rect 129834 301494 130454 334938
rect 129834 301258 129866 301494
rect 130102 301258 130186 301494
rect 130422 301258 130454 301494
rect 129834 301174 130454 301258
rect 129834 300938 129866 301174
rect 130102 300938 130186 301174
rect 130422 300938 130454 301174
rect 129834 267494 130454 300938
rect 129834 267258 129866 267494
rect 130102 267258 130186 267494
rect 130422 267258 130454 267494
rect 129834 267174 130454 267258
rect 129834 266938 129866 267174
rect 130102 266938 130186 267174
rect 130422 266938 130454 267174
rect 129834 233494 130454 266938
rect 129834 233258 129866 233494
rect 130102 233258 130186 233494
rect 130422 233258 130454 233494
rect 129834 233174 130454 233258
rect 129834 232938 129866 233174
rect 130102 232938 130186 233174
rect 130422 232938 130454 233174
rect 65300 225466 71300 225565
rect 43234 214658 43266 214894
rect 43502 214658 43586 214894
rect 43822 214658 43854 214894
rect 43234 214574 43854 214658
rect 43234 214338 43266 214574
rect 43502 214338 43586 214574
rect 43822 214338 43854 214574
rect 43234 180894 43854 214338
rect 43234 180658 43266 180894
rect 43502 180658 43586 180894
rect 43822 180658 43854 180894
rect 43234 180574 43854 180658
rect 43234 180338 43266 180574
rect 43502 180338 43586 180574
rect 43822 180338 43854 180574
rect 43234 146894 43854 180338
rect 43234 146658 43266 146894
rect 43502 146658 43586 146894
rect 43822 146658 43854 146894
rect 43234 146574 43854 146658
rect 43234 146338 43266 146574
rect 43502 146338 43586 146574
rect 43822 146338 43854 146574
rect 43234 112894 43854 146338
rect 43234 112658 43266 112894
rect 43502 112658 43586 112894
rect 43822 112658 43854 112894
rect 43234 112574 43854 112658
rect 43234 112338 43266 112574
rect 43502 112338 43586 112574
rect 43822 112338 43854 112574
rect 43234 78894 43854 112338
rect 43234 78658 43266 78894
rect 43502 78658 43586 78894
rect 43822 78658 43854 78894
rect 43234 78574 43854 78658
rect 43234 78338 43266 78574
rect 43502 78338 43586 78574
rect 43822 78338 43854 78574
rect 43234 44894 43854 78338
rect 43234 44658 43266 44894
rect 43502 44658 43586 44894
rect 43822 44658 43854 44894
rect 43234 44574 43854 44658
rect 43234 44338 43266 44574
rect 43502 44338 43586 44574
rect 43822 44338 43854 44574
rect 43234 10894 43854 44338
rect 43234 10658 43266 10894
rect 43502 10658 43586 10894
rect 43822 10658 43854 10894
rect 43234 10574 43854 10658
rect 43234 10338 43266 10574
rect 43502 10338 43586 10574
rect 43822 10338 43854 10574
rect 43234 -2266 43854 10338
rect 43234 -2502 43266 -2266
rect 43502 -2502 43586 -2266
rect 43822 -2502 43854 -2266
rect 43234 -2586 43854 -2502
rect 43234 -2822 43266 -2586
rect 43502 -2822 43586 -2586
rect 43822 -2822 43854 -2586
rect 43234 -7654 43854 -2822
rect 46954 184614 47574 214340
rect 46954 184378 46986 184614
rect 47222 184378 47306 184614
rect 47542 184378 47574 184614
rect 46954 184294 47574 184378
rect 46954 184058 46986 184294
rect 47222 184058 47306 184294
rect 47542 184058 47574 184294
rect 46954 150614 47574 184058
rect 46954 150378 46986 150614
rect 47222 150378 47306 150614
rect 47542 150378 47574 150614
rect 46954 150294 47574 150378
rect 46954 150058 46986 150294
rect 47222 150058 47306 150294
rect 47542 150058 47574 150294
rect 46954 116614 47574 150058
rect 46954 116378 46986 116614
rect 47222 116378 47306 116614
rect 47542 116378 47574 116614
rect 46954 116294 47574 116378
rect 46954 116058 46986 116294
rect 47222 116058 47306 116294
rect 47542 116058 47574 116294
rect 46954 82614 47574 116058
rect 46954 82378 46986 82614
rect 47222 82378 47306 82614
rect 47542 82378 47574 82614
rect 46954 82294 47574 82378
rect 46954 82058 46986 82294
rect 47222 82058 47306 82294
rect 47542 82058 47574 82294
rect 46954 48614 47574 82058
rect 46954 48378 46986 48614
rect 47222 48378 47306 48614
rect 47542 48378 47574 48614
rect 46954 48294 47574 48378
rect 46954 48058 46986 48294
rect 47222 48058 47306 48294
rect 47542 48058 47574 48294
rect 46954 14614 47574 48058
rect 46954 14378 46986 14614
rect 47222 14378 47306 14614
rect 47542 14378 47574 14614
rect 46954 14294 47574 14378
rect 46954 14058 46986 14294
rect 47222 14058 47306 14294
rect 47542 14058 47574 14294
rect 46954 -3226 47574 14058
rect 46954 -3462 46986 -3226
rect 47222 -3462 47306 -3226
rect 47542 -3462 47574 -3226
rect 46954 -3546 47574 -3462
rect 46954 -3782 46986 -3546
rect 47222 -3782 47306 -3546
rect 47542 -3782 47574 -3546
rect 46954 -7654 47574 -3782
rect 50674 188334 51294 214340
rect 50674 188098 50706 188334
rect 50942 188098 51026 188334
rect 51262 188098 51294 188334
rect 50674 188014 51294 188098
rect 50674 187778 50706 188014
rect 50942 187778 51026 188014
rect 51262 187778 51294 188014
rect 50674 154334 51294 187778
rect 50674 154098 50706 154334
rect 50942 154098 51026 154334
rect 51262 154098 51294 154334
rect 50674 154014 51294 154098
rect 50674 153778 50706 154014
rect 50942 153778 51026 154014
rect 51262 153778 51294 154014
rect 50674 120334 51294 153778
rect 50674 120098 50706 120334
rect 50942 120098 51026 120334
rect 51262 120098 51294 120334
rect 50674 120014 51294 120098
rect 50674 119778 50706 120014
rect 50942 119778 51026 120014
rect 51262 119778 51294 120014
rect 50674 86334 51294 119778
rect 50674 86098 50706 86334
rect 50942 86098 51026 86334
rect 51262 86098 51294 86334
rect 50674 86014 51294 86098
rect 50674 85778 50706 86014
rect 50942 85778 51026 86014
rect 51262 85778 51294 86014
rect 50674 52334 51294 85778
rect 50674 52098 50706 52334
rect 50942 52098 51026 52334
rect 51262 52098 51294 52334
rect 50674 52014 51294 52098
rect 50674 51778 50706 52014
rect 50942 51778 51026 52014
rect 51262 51778 51294 52014
rect 50674 18334 51294 51778
rect 50674 18098 50706 18334
rect 50942 18098 51026 18334
rect 51262 18098 51294 18334
rect 50674 18014 51294 18098
rect 50674 17778 50706 18014
rect 50942 17778 51026 18014
rect 51262 17778 51294 18014
rect 50674 -4186 51294 17778
rect 50674 -4422 50706 -4186
rect 50942 -4422 51026 -4186
rect 51262 -4422 51294 -4186
rect 50674 -4506 51294 -4422
rect 50674 -4742 50706 -4506
rect 50942 -4742 51026 -4506
rect 51262 -4742 51294 -4506
rect 50674 -7654 51294 -4742
rect 54394 192054 55014 214340
rect 54394 191818 54426 192054
rect 54662 191818 54746 192054
rect 54982 191818 55014 192054
rect 54394 191734 55014 191818
rect 54394 191498 54426 191734
rect 54662 191498 54746 191734
rect 54982 191498 55014 191734
rect 54394 158054 55014 191498
rect 54394 157818 54426 158054
rect 54662 157818 54746 158054
rect 54982 157818 55014 158054
rect 54394 157734 55014 157818
rect 54394 157498 54426 157734
rect 54662 157498 54746 157734
rect 54982 157498 55014 157734
rect 54394 124054 55014 157498
rect 54394 123818 54426 124054
rect 54662 123818 54746 124054
rect 54982 123818 55014 124054
rect 54394 123734 55014 123818
rect 54394 123498 54426 123734
rect 54662 123498 54746 123734
rect 54982 123498 55014 123734
rect 54394 90054 55014 123498
rect 54394 89818 54426 90054
rect 54662 89818 54746 90054
rect 54982 89818 55014 90054
rect 54394 89734 55014 89818
rect 54394 89498 54426 89734
rect 54662 89498 54746 89734
rect 54982 89498 55014 89734
rect 54394 56054 55014 89498
rect 54394 55818 54426 56054
rect 54662 55818 54746 56054
rect 54982 55818 55014 56054
rect 54394 55734 55014 55818
rect 54394 55498 54426 55734
rect 54662 55498 54746 55734
rect 54982 55498 55014 55734
rect 54394 22054 55014 55498
rect 54394 21818 54426 22054
rect 54662 21818 54746 22054
rect 54982 21818 55014 22054
rect 54394 21734 55014 21818
rect 54394 21498 54426 21734
rect 54662 21498 54746 21734
rect 54982 21498 55014 21734
rect 54394 -5146 55014 21498
rect 54394 -5382 54426 -5146
rect 54662 -5382 54746 -5146
rect 54982 -5382 55014 -5146
rect 54394 -5466 55014 -5382
rect 54394 -5702 54426 -5466
rect 54662 -5702 54746 -5466
rect 54982 -5702 55014 -5466
rect 54394 -7654 55014 -5702
rect 58114 195774 58734 214340
rect 58114 195538 58146 195774
rect 58382 195538 58466 195774
rect 58702 195538 58734 195774
rect 58114 195454 58734 195538
rect 58114 195218 58146 195454
rect 58382 195218 58466 195454
rect 58702 195218 58734 195454
rect 58114 161774 58734 195218
rect 58114 161538 58146 161774
rect 58382 161538 58466 161774
rect 58702 161538 58734 161774
rect 58114 161454 58734 161538
rect 58114 161218 58146 161454
rect 58382 161218 58466 161454
rect 58702 161218 58734 161454
rect 58114 127774 58734 161218
rect 58114 127538 58146 127774
rect 58382 127538 58466 127774
rect 58702 127538 58734 127774
rect 58114 127454 58734 127538
rect 58114 127218 58146 127454
rect 58382 127218 58466 127454
rect 58702 127218 58734 127454
rect 58114 93774 58734 127218
rect 58114 93538 58146 93774
rect 58382 93538 58466 93774
rect 58702 93538 58734 93774
rect 58114 93454 58734 93538
rect 58114 93218 58146 93454
rect 58382 93218 58466 93454
rect 58702 93218 58734 93454
rect 58114 59774 58734 93218
rect 58114 59538 58146 59774
rect 58382 59538 58466 59774
rect 58702 59538 58734 59774
rect 58114 59454 58734 59538
rect 58114 59218 58146 59454
rect 58382 59218 58466 59454
rect 58702 59218 58734 59454
rect 58114 25774 58734 59218
rect 58114 25538 58146 25774
rect 58382 25538 58466 25774
rect 58702 25538 58734 25774
rect 58114 25454 58734 25538
rect 58114 25218 58146 25454
rect 58382 25218 58466 25454
rect 58702 25218 58734 25454
rect 58114 -6106 58734 25218
rect 58114 -6342 58146 -6106
rect 58382 -6342 58466 -6106
rect 58702 -6342 58734 -6106
rect 58114 -6426 58734 -6342
rect 58114 -6662 58146 -6426
rect 58382 -6662 58466 -6426
rect 58702 -6662 58734 -6426
rect 58114 -7654 58734 -6662
rect 61834 199494 62454 214340
rect 61834 199258 61866 199494
rect 62102 199258 62186 199494
rect 62422 199258 62454 199494
rect 61834 199174 62454 199258
rect 61834 198938 61866 199174
rect 62102 198938 62186 199174
rect 62422 198938 62454 199174
rect 61834 165494 62454 198938
rect 61834 165258 61866 165494
rect 62102 165258 62186 165494
rect 62422 165258 62454 165494
rect 61834 165174 62454 165258
rect 61834 164938 61866 165174
rect 62102 164938 62186 165174
rect 62422 164938 62454 165174
rect 61834 131494 62454 164938
rect 61834 131258 61866 131494
rect 62102 131258 62186 131494
rect 62422 131258 62454 131494
rect 61834 131174 62454 131258
rect 61834 130938 61866 131174
rect 62102 130938 62186 131174
rect 62422 130938 62454 131174
rect 61834 97494 62454 130938
rect 61834 97258 61866 97494
rect 62102 97258 62186 97494
rect 62422 97258 62454 97494
rect 61834 97174 62454 97258
rect 61834 96938 61866 97174
rect 62102 96938 62186 97174
rect 62422 96938 62454 97174
rect 61834 63494 62454 96938
rect 61834 63258 61866 63494
rect 62102 63258 62186 63494
rect 62422 63258 62454 63494
rect 61834 63174 62454 63258
rect 61834 62938 61866 63174
rect 62102 62938 62186 63174
rect 62422 62938 62454 63174
rect 61834 29494 62454 62938
rect 61834 29258 61866 29494
rect 62102 29258 62186 29494
rect 62422 29258 62454 29494
rect 61834 29174 62454 29258
rect 61834 28938 61866 29174
rect 62102 28938 62186 29174
rect 62422 28938 62454 29174
rect 61834 -7066 62454 28938
rect 61834 -7302 61866 -7066
rect 62102 -7302 62186 -7066
rect 62422 -7302 62454 -7066
rect 61834 -7386 62454 -7302
rect 61834 -7622 61866 -7386
rect 62102 -7622 62186 -7386
rect 62422 -7622 62454 -7386
rect 61834 -7654 62454 -7622
rect 69794 207454 70414 223020
rect 69794 207218 69826 207454
rect 70062 207218 70146 207454
rect 70382 207218 70414 207454
rect 69794 207134 70414 207218
rect 69794 206898 69826 207134
rect 70062 206898 70146 207134
rect 70382 206898 70414 207134
rect 69794 173454 70414 206898
rect 69794 173218 69826 173454
rect 70062 173218 70146 173454
rect 70382 173218 70414 173454
rect 69794 173134 70414 173218
rect 69794 172898 69826 173134
rect 70062 172898 70146 173134
rect 70382 172898 70414 173134
rect 69794 139454 70414 172898
rect 69794 139218 69826 139454
rect 70062 139218 70146 139454
rect 70382 139218 70414 139454
rect 69794 139134 70414 139218
rect 69794 138898 69826 139134
rect 70062 138898 70146 139134
rect 70382 138898 70414 139134
rect 69794 105454 70414 138898
rect 69794 105218 69826 105454
rect 70062 105218 70146 105454
rect 70382 105218 70414 105454
rect 69794 105134 70414 105218
rect 69794 104898 69826 105134
rect 70062 104898 70146 105134
rect 70382 104898 70414 105134
rect 69794 71454 70414 104898
rect 69794 71218 69826 71454
rect 70062 71218 70146 71454
rect 70382 71218 70414 71454
rect 69794 71134 70414 71218
rect 69794 70898 69826 71134
rect 70062 70898 70146 71134
rect 70382 70898 70414 71134
rect 69794 37454 70414 70898
rect 69794 37218 69826 37454
rect 70062 37218 70146 37454
rect 70382 37218 70414 37454
rect 69794 37134 70414 37218
rect 69794 36898 69826 37134
rect 70062 36898 70146 37134
rect 70382 36898 70414 37134
rect 69794 3454 70414 36898
rect 69794 3218 69826 3454
rect 70062 3218 70146 3454
rect 70382 3218 70414 3454
rect 69794 3134 70414 3218
rect 69794 2898 69826 3134
rect 70062 2898 70146 3134
rect 70382 2898 70414 3134
rect 69794 -346 70414 2898
rect 69794 -582 69826 -346
rect 70062 -582 70146 -346
rect 70382 -582 70414 -346
rect 69794 -666 70414 -582
rect 69794 -902 69826 -666
rect 70062 -902 70146 -666
rect 70382 -902 70414 -666
rect 69794 -7654 70414 -902
rect 73514 211174 74134 214340
rect 73514 210938 73546 211174
rect 73782 210938 73866 211174
rect 74102 210938 74134 211174
rect 73514 210854 74134 210938
rect 73514 210618 73546 210854
rect 73782 210618 73866 210854
rect 74102 210618 74134 210854
rect 73514 177174 74134 210618
rect 73514 176938 73546 177174
rect 73782 176938 73866 177174
rect 74102 176938 74134 177174
rect 73514 176854 74134 176938
rect 73514 176618 73546 176854
rect 73782 176618 73866 176854
rect 74102 176618 74134 176854
rect 73514 143174 74134 176618
rect 73514 142938 73546 143174
rect 73782 142938 73866 143174
rect 74102 142938 74134 143174
rect 73514 142854 74134 142938
rect 73514 142618 73546 142854
rect 73782 142618 73866 142854
rect 74102 142618 74134 142854
rect 73514 109174 74134 142618
rect 73514 108938 73546 109174
rect 73782 108938 73866 109174
rect 74102 108938 74134 109174
rect 73514 108854 74134 108938
rect 73514 108618 73546 108854
rect 73782 108618 73866 108854
rect 74102 108618 74134 108854
rect 73514 75174 74134 108618
rect 73514 74938 73546 75174
rect 73782 74938 73866 75174
rect 74102 74938 74134 75174
rect 73514 74854 74134 74938
rect 73514 74618 73546 74854
rect 73782 74618 73866 74854
rect 74102 74618 74134 74854
rect 73514 41174 74134 74618
rect 73514 40938 73546 41174
rect 73782 40938 73866 41174
rect 74102 40938 74134 41174
rect 73514 40854 74134 40938
rect 73514 40618 73546 40854
rect 73782 40618 73866 40854
rect 74102 40618 74134 40854
rect 73514 7174 74134 40618
rect 73514 6938 73546 7174
rect 73782 6938 73866 7174
rect 74102 6938 74134 7174
rect 73514 6854 74134 6938
rect 73514 6618 73546 6854
rect 73782 6618 73866 6854
rect 74102 6618 74134 6854
rect 73514 -1306 74134 6618
rect 73514 -1542 73546 -1306
rect 73782 -1542 73866 -1306
rect 74102 -1542 74134 -1306
rect 73514 -1626 74134 -1542
rect 73514 -1862 73546 -1626
rect 73782 -1862 73866 -1626
rect 74102 -1862 74134 -1626
rect 73514 -7654 74134 -1862
rect 77234 180894 77854 214340
rect 77234 180658 77266 180894
rect 77502 180658 77586 180894
rect 77822 180658 77854 180894
rect 77234 180574 77854 180658
rect 77234 180338 77266 180574
rect 77502 180338 77586 180574
rect 77822 180338 77854 180574
rect 77234 146894 77854 180338
rect 77234 146658 77266 146894
rect 77502 146658 77586 146894
rect 77822 146658 77854 146894
rect 77234 146574 77854 146658
rect 77234 146338 77266 146574
rect 77502 146338 77586 146574
rect 77822 146338 77854 146574
rect 77234 112894 77854 146338
rect 77234 112658 77266 112894
rect 77502 112658 77586 112894
rect 77822 112658 77854 112894
rect 77234 112574 77854 112658
rect 77234 112338 77266 112574
rect 77502 112338 77586 112574
rect 77822 112338 77854 112574
rect 77234 78894 77854 112338
rect 77234 78658 77266 78894
rect 77502 78658 77586 78894
rect 77822 78658 77854 78894
rect 77234 78574 77854 78658
rect 77234 78338 77266 78574
rect 77502 78338 77586 78574
rect 77822 78338 77854 78574
rect 77234 44894 77854 78338
rect 77234 44658 77266 44894
rect 77502 44658 77586 44894
rect 77822 44658 77854 44894
rect 77234 44574 77854 44658
rect 77234 44338 77266 44574
rect 77502 44338 77586 44574
rect 77822 44338 77854 44574
rect 77234 10894 77854 44338
rect 77234 10658 77266 10894
rect 77502 10658 77586 10894
rect 77822 10658 77854 10894
rect 77234 10574 77854 10658
rect 77234 10338 77266 10574
rect 77502 10338 77586 10574
rect 77822 10338 77854 10574
rect 77234 -2266 77854 10338
rect 77234 -2502 77266 -2266
rect 77502 -2502 77586 -2266
rect 77822 -2502 77854 -2266
rect 77234 -2586 77854 -2502
rect 77234 -2822 77266 -2586
rect 77502 -2822 77586 -2586
rect 77822 -2822 77854 -2586
rect 77234 -7654 77854 -2822
rect 80954 184614 81574 214340
rect 80954 184378 80986 184614
rect 81222 184378 81306 184614
rect 81542 184378 81574 184614
rect 80954 184294 81574 184378
rect 80954 184058 80986 184294
rect 81222 184058 81306 184294
rect 81542 184058 81574 184294
rect 80954 150614 81574 184058
rect 80954 150378 80986 150614
rect 81222 150378 81306 150614
rect 81542 150378 81574 150614
rect 80954 150294 81574 150378
rect 80954 150058 80986 150294
rect 81222 150058 81306 150294
rect 81542 150058 81574 150294
rect 80954 116614 81574 150058
rect 80954 116378 80986 116614
rect 81222 116378 81306 116614
rect 81542 116378 81574 116614
rect 80954 116294 81574 116378
rect 80954 116058 80986 116294
rect 81222 116058 81306 116294
rect 81542 116058 81574 116294
rect 80954 82614 81574 116058
rect 80954 82378 80986 82614
rect 81222 82378 81306 82614
rect 81542 82378 81574 82614
rect 80954 82294 81574 82378
rect 80954 82058 80986 82294
rect 81222 82058 81306 82294
rect 81542 82058 81574 82294
rect 80954 48614 81574 82058
rect 80954 48378 80986 48614
rect 81222 48378 81306 48614
rect 81542 48378 81574 48614
rect 80954 48294 81574 48378
rect 80954 48058 80986 48294
rect 81222 48058 81306 48294
rect 81542 48058 81574 48294
rect 80954 14614 81574 48058
rect 80954 14378 80986 14614
rect 81222 14378 81306 14614
rect 81542 14378 81574 14614
rect 80954 14294 81574 14378
rect 80954 14058 80986 14294
rect 81222 14058 81306 14294
rect 81542 14058 81574 14294
rect 80954 -3226 81574 14058
rect 80954 -3462 80986 -3226
rect 81222 -3462 81306 -3226
rect 81542 -3462 81574 -3226
rect 80954 -3546 81574 -3462
rect 80954 -3782 80986 -3546
rect 81222 -3782 81306 -3546
rect 81542 -3782 81574 -3546
rect 80954 -7654 81574 -3782
rect 84674 188334 85294 214340
rect 84674 188098 84706 188334
rect 84942 188098 85026 188334
rect 85262 188098 85294 188334
rect 84674 188014 85294 188098
rect 84674 187778 84706 188014
rect 84942 187778 85026 188014
rect 85262 187778 85294 188014
rect 84674 154334 85294 187778
rect 84674 154098 84706 154334
rect 84942 154098 85026 154334
rect 85262 154098 85294 154334
rect 84674 154014 85294 154098
rect 84674 153778 84706 154014
rect 84942 153778 85026 154014
rect 85262 153778 85294 154014
rect 84674 120334 85294 153778
rect 84674 120098 84706 120334
rect 84942 120098 85026 120334
rect 85262 120098 85294 120334
rect 84674 120014 85294 120098
rect 84674 119778 84706 120014
rect 84942 119778 85026 120014
rect 85262 119778 85294 120014
rect 84674 86334 85294 119778
rect 84674 86098 84706 86334
rect 84942 86098 85026 86334
rect 85262 86098 85294 86334
rect 84674 86014 85294 86098
rect 84674 85778 84706 86014
rect 84942 85778 85026 86014
rect 85262 85778 85294 86014
rect 84674 52334 85294 85778
rect 84674 52098 84706 52334
rect 84942 52098 85026 52334
rect 85262 52098 85294 52334
rect 84674 52014 85294 52098
rect 84674 51778 84706 52014
rect 84942 51778 85026 52014
rect 85262 51778 85294 52014
rect 84674 18334 85294 51778
rect 84674 18098 84706 18334
rect 84942 18098 85026 18334
rect 85262 18098 85294 18334
rect 84674 18014 85294 18098
rect 84674 17778 84706 18014
rect 84942 17778 85026 18014
rect 85262 17778 85294 18014
rect 84674 -4186 85294 17778
rect 84674 -4422 84706 -4186
rect 84942 -4422 85026 -4186
rect 85262 -4422 85294 -4186
rect 84674 -4506 85294 -4422
rect 84674 -4742 84706 -4506
rect 84942 -4742 85026 -4506
rect 85262 -4742 85294 -4506
rect 84674 -7654 85294 -4742
rect 88394 192054 89014 214340
rect 88394 191818 88426 192054
rect 88662 191818 88746 192054
rect 88982 191818 89014 192054
rect 88394 191734 89014 191818
rect 88394 191498 88426 191734
rect 88662 191498 88746 191734
rect 88982 191498 89014 191734
rect 88394 158054 89014 191498
rect 88394 157818 88426 158054
rect 88662 157818 88746 158054
rect 88982 157818 89014 158054
rect 88394 157734 89014 157818
rect 88394 157498 88426 157734
rect 88662 157498 88746 157734
rect 88982 157498 89014 157734
rect 88394 124054 89014 157498
rect 88394 123818 88426 124054
rect 88662 123818 88746 124054
rect 88982 123818 89014 124054
rect 88394 123734 89014 123818
rect 88394 123498 88426 123734
rect 88662 123498 88746 123734
rect 88982 123498 89014 123734
rect 88394 90054 89014 123498
rect 88394 89818 88426 90054
rect 88662 89818 88746 90054
rect 88982 89818 89014 90054
rect 88394 89734 89014 89818
rect 88394 89498 88426 89734
rect 88662 89498 88746 89734
rect 88982 89498 89014 89734
rect 88394 56054 89014 89498
rect 88394 55818 88426 56054
rect 88662 55818 88746 56054
rect 88982 55818 89014 56054
rect 88394 55734 89014 55818
rect 88394 55498 88426 55734
rect 88662 55498 88746 55734
rect 88982 55498 89014 55734
rect 88394 22054 89014 55498
rect 88394 21818 88426 22054
rect 88662 21818 88746 22054
rect 88982 21818 89014 22054
rect 88394 21734 89014 21818
rect 88394 21498 88426 21734
rect 88662 21498 88746 21734
rect 88982 21498 89014 21734
rect 88394 -5146 89014 21498
rect 88394 -5382 88426 -5146
rect 88662 -5382 88746 -5146
rect 88982 -5382 89014 -5146
rect 88394 -5466 89014 -5382
rect 88394 -5702 88426 -5466
rect 88662 -5702 88746 -5466
rect 88982 -5702 89014 -5466
rect 88394 -7654 89014 -5702
rect 92114 195774 92734 214340
rect 92114 195538 92146 195774
rect 92382 195538 92466 195774
rect 92702 195538 92734 195774
rect 92114 195454 92734 195538
rect 92114 195218 92146 195454
rect 92382 195218 92466 195454
rect 92702 195218 92734 195454
rect 92114 161774 92734 195218
rect 92114 161538 92146 161774
rect 92382 161538 92466 161774
rect 92702 161538 92734 161774
rect 92114 161454 92734 161538
rect 92114 161218 92146 161454
rect 92382 161218 92466 161454
rect 92702 161218 92734 161454
rect 92114 127774 92734 161218
rect 92114 127538 92146 127774
rect 92382 127538 92466 127774
rect 92702 127538 92734 127774
rect 92114 127454 92734 127538
rect 92114 127218 92146 127454
rect 92382 127218 92466 127454
rect 92702 127218 92734 127454
rect 92114 93774 92734 127218
rect 92114 93538 92146 93774
rect 92382 93538 92466 93774
rect 92702 93538 92734 93774
rect 92114 93454 92734 93538
rect 92114 93218 92146 93454
rect 92382 93218 92466 93454
rect 92702 93218 92734 93454
rect 92114 59774 92734 93218
rect 92114 59538 92146 59774
rect 92382 59538 92466 59774
rect 92702 59538 92734 59774
rect 92114 59454 92734 59538
rect 92114 59218 92146 59454
rect 92382 59218 92466 59454
rect 92702 59218 92734 59454
rect 92114 25774 92734 59218
rect 92114 25538 92146 25774
rect 92382 25538 92466 25774
rect 92702 25538 92734 25774
rect 92114 25454 92734 25538
rect 92114 25218 92146 25454
rect 92382 25218 92466 25454
rect 92702 25218 92734 25454
rect 92114 -6106 92734 25218
rect 92114 -6342 92146 -6106
rect 92382 -6342 92466 -6106
rect 92702 -6342 92734 -6106
rect 92114 -6426 92734 -6342
rect 92114 -6662 92146 -6426
rect 92382 -6662 92466 -6426
rect 92702 -6662 92734 -6426
rect 92114 -7654 92734 -6662
rect 95834 199494 96454 214340
rect 95834 199258 95866 199494
rect 96102 199258 96186 199494
rect 96422 199258 96454 199494
rect 95834 199174 96454 199258
rect 95834 198938 95866 199174
rect 96102 198938 96186 199174
rect 96422 198938 96454 199174
rect 95834 165494 96454 198938
rect 95834 165258 95866 165494
rect 96102 165258 96186 165494
rect 96422 165258 96454 165494
rect 95834 165174 96454 165258
rect 95834 164938 95866 165174
rect 96102 164938 96186 165174
rect 96422 164938 96454 165174
rect 95834 131494 96454 164938
rect 95834 131258 95866 131494
rect 96102 131258 96186 131494
rect 96422 131258 96454 131494
rect 95834 131174 96454 131258
rect 95834 130938 95866 131174
rect 96102 130938 96186 131174
rect 96422 130938 96454 131174
rect 95834 97494 96454 130938
rect 95834 97258 95866 97494
rect 96102 97258 96186 97494
rect 96422 97258 96454 97494
rect 95834 97174 96454 97258
rect 95834 96938 95866 97174
rect 96102 96938 96186 97174
rect 96422 96938 96454 97174
rect 95834 63494 96454 96938
rect 95834 63258 95866 63494
rect 96102 63258 96186 63494
rect 96422 63258 96454 63494
rect 95834 63174 96454 63258
rect 95834 62938 95866 63174
rect 96102 62938 96186 63174
rect 96422 62938 96454 63174
rect 95834 29494 96454 62938
rect 95834 29258 95866 29494
rect 96102 29258 96186 29494
rect 96422 29258 96454 29494
rect 95834 29174 96454 29258
rect 95834 28938 95866 29174
rect 96102 28938 96186 29174
rect 96422 28938 96454 29174
rect 95834 -7066 96454 28938
rect 95834 -7302 95866 -7066
rect 96102 -7302 96186 -7066
rect 96422 -7302 96454 -7066
rect 95834 -7386 96454 -7302
rect 95834 -7622 95866 -7386
rect 96102 -7622 96186 -7386
rect 96422 -7622 96454 -7386
rect 95834 -7654 96454 -7622
rect 103794 207454 104414 214340
rect 103794 207218 103826 207454
rect 104062 207218 104146 207454
rect 104382 207218 104414 207454
rect 103794 207134 104414 207218
rect 103794 206898 103826 207134
rect 104062 206898 104146 207134
rect 104382 206898 104414 207134
rect 103794 173454 104414 206898
rect 103794 173218 103826 173454
rect 104062 173218 104146 173454
rect 104382 173218 104414 173454
rect 103794 173134 104414 173218
rect 103794 172898 103826 173134
rect 104062 172898 104146 173134
rect 104382 172898 104414 173134
rect 103794 139454 104414 172898
rect 103794 139218 103826 139454
rect 104062 139218 104146 139454
rect 104382 139218 104414 139454
rect 103794 139134 104414 139218
rect 103794 138898 103826 139134
rect 104062 138898 104146 139134
rect 104382 138898 104414 139134
rect 103794 105454 104414 138898
rect 103794 105218 103826 105454
rect 104062 105218 104146 105454
rect 104382 105218 104414 105454
rect 103794 105134 104414 105218
rect 103794 104898 103826 105134
rect 104062 104898 104146 105134
rect 104382 104898 104414 105134
rect 103794 71454 104414 104898
rect 103794 71218 103826 71454
rect 104062 71218 104146 71454
rect 104382 71218 104414 71454
rect 103794 71134 104414 71218
rect 103794 70898 103826 71134
rect 104062 70898 104146 71134
rect 104382 70898 104414 71134
rect 103794 37454 104414 70898
rect 103794 37218 103826 37454
rect 104062 37218 104146 37454
rect 104382 37218 104414 37454
rect 103794 37134 104414 37218
rect 103794 36898 103826 37134
rect 104062 36898 104146 37134
rect 104382 36898 104414 37134
rect 103794 3454 104414 36898
rect 103794 3218 103826 3454
rect 104062 3218 104146 3454
rect 104382 3218 104414 3454
rect 103794 3134 104414 3218
rect 103794 2898 103826 3134
rect 104062 2898 104146 3134
rect 104382 2898 104414 3134
rect 103794 -346 104414 2898
rect 103794 -582 103826 -346
rect 104062 -582 104146 -346
rect 104382 -582 104414 -346
rect 103794 -666 104414 -582
rect 103794 -902 103826 -666
rect 104062 -902 104146 -666
rect 104382 -902 104414 -666
rect 103794 -7654 104414 -902
rect 107514 211174 108134 214340
rect 107514 210938 107546 211174
rect 107782 210938 107866 211174
rect 108102 210938 108134 211174
rect 107514 210854 108134 210938
rect 107514 210618 107546 210854
rect 107782 210618 107866 210854
rect 108102 210618 108134 210854
rect 107514 177174 108134 210618
rect 107514 176938 107546 177174
rect 107782 176938 107866 177174
rect 108102 176938 108134 177174
rect 107514 176854 108134 176938
rect 107514 176618 107546 176854
rect 107782 176618 107866 176854
rect 108102 176618 108134 176854
rect 107514 143174 108134 176618
rect 107514 142938 107546 143174
rect 107782 142938 107866 143174
rect 108102 142938 108134 143174
rect 107514 142854 108134 142938
rect 107514 142618 107546 142854
rect 107782 142618 107866 142854
rect 108102 142618 108134 142854
rect 107514 109174 108134 142618
rect 107514 108938 107546 109174
rect 107782 108938 107866 109174
rect 108102 108938 108134 109174
rect 107514 108854 108134 108938
rect 107514 108618 107546 108854
rect 107782 108618 107866 108854
rect 108102 108618 108134 108854
rect 107514 75174 108134 108618
rect 107514 74938 107546 75174
rect 107782 74938 107866 75174
rect 108102 74938 108134 75174
rect 107514 74854 108134 74938
rect 107514 74618 107546 74854
rect 107782 74618 107866 74854
rect 108102 74618 108134 74854
rect 107514 41174 108134 74618
rect 107514 40938 107546 41174
rect 107782 40938 107866 41174
rect 108102 40938 108134 41174
rect 107514 40854 108134 40938
rect 107514 40618 107546 40854
rect 107782 40618 107866 40854
rect 108102 40618 108134 40854
rect 107514 7174 108134 40618
rect 107514 6938 107546 7174
rect 107782 6938 107866 7174
rect 108102 6938 108134 7174
rect 107514 6854 108134 6938
rect 107514 6618 107546 6854
rect 107782 6618 107866 6854
rect 108102 6618 108134 6854
rect 107514 -1306 108134 6618
rect 107514 -1542 107546 -1306
rect 107782 -1542 107866 -1306
rect 108102 -1542 108134 -1306
rect 107514 -1626 108134 -1542
rect 107514 -1862 107546 -1626
rect 107782 -1862 107866 -1626
rect 108102 -1862 108134 -1626
rect 107514 -7654 108134 -1862
rect 111234 180894 111854 214340
rect 111234 180658 111266 180894
rect 111502 180658 111586 180894
rect 111822 180658 111854 180894
rect 111234 180574 111854 180658
rect 111234 180338 111266 180574
rect 111502 180338 111586 180574
rect 111822 180338 111854 180574
rect 111234 146894 111854 180338
rect 111234 146658 111266 146894
rect 111502 146658 111586 146894
rect 111822 146658 111854 146894
rect 111234 146574 111854 146658
rect 111234 146338 111266 146574
rect 111502 146338 111586 146574
rect 111822 146338 111854 146574
rect 111234 112894 111854 146338
rect 111234 112658 111266 112894
rect 111502 112658 111586 112894
rect 111822 112658 111854 112894
rect 111234 112574 111854 112658
rect 111234 112338 111266 112574
rect 111502 112338 111586 112574
rect 111822 112338 111854 112574
rect 111234 78894 111854 112338
rect 111234 78658 111266 78894
rect 111502 78658 111586 78894
rect 111822 78658 111854 78894
rect 111234 78574 111854 78658
rect 111234 78338 111266 78574
rect 111502 78338 111586 78574
rect 111822 78338 111854 78574
rect 111234 44894 111854 78338
rect 111234 44658 111266 44894
rect 111502 44658 111586 44894
rect 111822 44658 111854 44894
rect 111234 44574 111854 44658
rect 111234 44338 111266 44574
rect 111502 44338 111586 44574
rect 111822 44338 111854 44574
rect 111234 10894 111854 44338
rect 111234 10658 111266 10894
rect 111502 10658 111586 10894
rect 111822 10658 111854 10894
rect 111234 10574 111854 10658
rect 111234 10338 111266 10574
rect 111502 10338 111586 10574
rect 111822 10338 111854 10574
rect 111234 -2266 111854 10338
rect 111234 -2502 111266 -2266
rect 111502 -2502 111586 -2266
rect 111822 -2502 111854 -2266
rect 111234 -2586 111854 -2502
rect 111234 -2822 111266 -2586
rect 111502 -2822 111586 -2586
rect 111822 -2822 111854 -2586
rect 111234 -7654 111854 -2822
rect 114954 184614 115574 214340
rect 114954 184378 114986 184614
rect 115222 184378 115306 184614
rect 115542 184378 115574 184614
rect 114954 184294 115574 184378
rect 114954 184058 114986 184294
rect 115222 184058 115306 184294
rect 115542 184058 115574 184294
rect 114954 150614 115574 184058
rect 114954 150378 114986 150614
rect 115222 150378 115306 150614
rect 115542 150378 115574 150614
rect 114954 150294 115574 150378
rect 114954 150058 114986 150294
rect 115222 150058 115306 150294
rect 115542 150058 115574 150294
rect 114954 116614 115574 150058
rect 118674 188334 119294 214340
rect 118674 188098 118706 188334
rect 118942 188098 119026 188334
rect 119262 188098 119294 188334
rect 118674 188014 119294 188098
rect 118674 187778 118706 188014
rect 118942 187778 119026 188014
rect 119262 187778 119294 188014
rect 118674 154334 119294 187778
rect 118674 154098 118706 154334
rect 118942 154098 119026 154334
rect 119262 154098 119294 154334
rect 118674 154014 119294 154098
rect 118674 153778 118706 154014
rect 118942 153778 119026 154014
rect 119262 153778 119294 154014
rect 118674 134417 119294 153778
rect 122394 192054 123014 214340
rect 122394 191818 122426 192054
rect 122662 191818 122746 192054
rect 122982 191818 123014 192054
rect 122394 191734 123014 191818
rect 122394 191498 122426 191734
rect 122662 191498 122746 191734
rect 122982 191498 123014 191734
rect 122394 158054 123014 191498
rect 122394 157818 122426 158054
rect 122662 157818 122746 158054
rect 122982 157818 123014 158054
rect 122394 157734 123014 157818
rect 122394 157498 122426 157734
rect 122662 157498 122746 157734
rect 122982 157498 123014 157734
rect 122394 134417 123014 157498
rect 126114 195774 126734 214340
rect 126114 195538 126146 195774
rect 126382 195538 126466 195774
rect 126702 195538 126734 195774
rect 126114 195454 126734 195538
rect 126114 195218 126146 195454
rect 126382 195218 126466 195454
rect 126702 195218 126734 195454
rect 126114 161774 126734 195218
rect 126114 161538 126146 161774
rect 126382 161538 126466 161774
rect 126702 161538 126734 161774
rect 126114 161454 126734 161538
rect 126114 161218 126146 161454
rect 126382 161218 126466 161454
rect 126702 161218 126734 161454
rect 126114 134417 126734 161218
rect 129834 199494 130454 232938
rect 137794 704838 138414 711590
rect 137794 704602 137826 704838
rect 138062 704602 138146 704838
rect 138382 704602 138414 704838
rect 137794 704518 138414 704602
rect 137794 704282 137826 704518
rect 138062 704282 138146 704518
rect 138382 704282 138414 704518
rect 137794 683454 138414 704282
rect 137794 683218 137826 683454
rect 138062 683218 138146 683454
rect 138382 683218 138414 683454
rect 137794 683134 138414 683218
rect 137794 682898 137826 683134
rect 138062 682898 138146 683134
rect 138382 682898 138414 683134
rect 137794 649454 138414 682898
rect 137794 649218 137826 649454
rect 138062 649218 138146 649454
rect 138382 649218 138414 649454
rect 137794 649134 138414 649218
rect 137794 648898 137826 649134
rect 138062 648898 138146 649134
rect 138382 648898 138414 649134
rect 137794 615454 138414 648898
rect 137794 615218 137826 615454
rect 138062 615218 138146 615454
rect 138382 615218 138414 615454
rect 137794 615134 138414 615218
rect 137794 614898 137826 615134
rect 138062 614898 138146 615134
rect 138382 614898 138414 615134
rect 137794 581454 138414 614898
rect 137794 581218 137826 581454
rect 138062 581218 138146 581454
rect 138382 581218 138414 581454
rect 137794 581134 138414 581218
rect 137794 580898 137826 581134
rect 138062 580898 138146 581134
rect 138382 580898 138414 581134
rect 137794 547454 138414 580898
rect 137794 547218 137826 547454
rect 138062 547218 138146 547454
rect 138382 547218 138414 547454
rect 137794 547134 138414 547218
rect 137794 546898 137826 547134
rect 138062 546898 138146 547134
rect 138382 546898 138414 547134
rect 137794 513454 138414 546898
rect 137794 513218 137826 513454
rect 138062 513218 138146 513454
rect 138382 513218 138414 513454
rect 137794 513134 138414 513218
rect 137794 512898 137826 513134
rect 138062 512898 138146 513134
rect 138382 512898 138414 513134
rect 137794 479454 138414 512898
rect 137794 479218 137826 479454
rect 138062 479218 138146 479454
rect 138382 479218 138414 479454
rect 137794 479134 138414 479218
rect 137794 478898 137826 479134
rect 138062 478898 138146 479134
rect 138382 478898 138414 479134
rect 137794 445454 138414 478898
rect 137794 445218 137826 445454
rect 138062 445218 138146 445454
rect 138382 445218 138414 445454
rect 137794 445134 138414 445218
rect 137794 444898 137826 445134
rect 138062 444898 138146 445134
rect 138382 444898 138414 445134
rect 137794 411454 138414 444898
rect 137794 411218 137826 411454
rect 138062 411218 138146 411454
rect 138382 411218 138414 411454
rect 137794 411134 138414 411218
rect 137794 410898 137826 411134
rect 138062 410898 138146 411134
rect 138382 410898 138414 411134
rect 137794 377454 138414 410898
rect 137794 377218 137826 377454
rect 138062 377218 138146 377454
rect 138382 377218 138414 377454
rect 137794 377134 138414 377218
rect 137794 376898 137826 377134
rect 138062 376898 138146 377134
rect 138382 376898 138414 377134
rect 137794 343454 138414 376898
rect 137794 343218 137826 343454
rect 138062 343218 138146 343454
rect 138382 343218 138414 343454
rect 137794 343134 138414 343218
rect 137794 342898 137826 343134
rect 138062 342898 138146 343134
rect 138382 342898 138414 343134
rect 137794 309454 138414 342898
rect 137794 309218 137826 309454
rect 138062 309218 138146 309454
rect 138382 309218 138414 309454
rect 137794 309134 138414 309218
rect 137794 308898 137826 309134
rect 138062 308898 138146 309134
rect 138382 308898 138414 309134
rect 137794 275454 138414 308898
rect 137794 275218 137826 275454
rect 138062 275218 138146 275454
rect 138382 275218 138414 275454
rect 137794 275134 138414 275218
rect 137794 274898 137826 275134
rect 138062 274898 138146 275134
rect 138382 274898 138414 275134
rect 137794 241454 138414 274898
rect 137794 241218 137826 241454
rect 138062 241218 138146 241454
rect 138382 241218 138414 241454
rect 137794 241134 138414 241218
rect 137794 240898 137826 241134
rect 138062 240898 138146 241134
rect 138382 240898 138414 241134
rect 137794 225660 138414 240898
rect 141514 705798 142134 711590
rect 141514 705562 141546 705798
rect 141782 705562 141866 705798
rect 142102 705562 142134 705798
rect 141514 705478 142134 705562
rect 141514 705242 141546 705478
rect 141782 705242 141866 705478
rect 142102 705242 142134 705478
rect 141514 687174 142134 705242
rect 141514 686938 141546 687174
rect 141782 686938 141866 687174
rect 142102 686938 142134 687174
rect 141514 686854 142134 686938
rect 141514 686618 141546 686854
rect 141782 686618 141866 686854
rect 142102 686618 142134 686854
rect 141514 653174 142134 686618
rect 141514 652938 141546 653174
rect 141782 652938 141866 653174
rect 142102 652938 142134 653174
rect 141514 652854 142134 652938
rect 141514 652618 141546 652854
rect 141782 652618 141866 652854
rect 142102 652618 142134 652854
rect 141514 619174 142134 652618
rect 141514 618938 141546 619174
rect 141782 618938 141866 619174
rect 142102 618938 142134 619174
rect 141514 618854 142134 618938
rect 141514 618618 141546 618854
rect 141782 618618 141866 618854
rect 142102 618618 142134 618854
rect 141514 585174 142134 618618
rect 141514 584938 141546 585174
rect 141782 584938 141866 585174
rect 142102 584938 142134 585174
rect 141514 584854 142134 584938
rect 141514 584618 141546 584854
rect 141782 584618 141866 584854
rect 142102 584618 142134 584854
rect 141514 551174 142134 584618
rect 141514 550938 141546 551174
rect 141782 550938 141866 551174
rect 142102 550938 142134 551174
rect 141514 550854 142134 550938
rect 141514 550618 141546 550854
rect 141782 550618 141866 550854
rect 142102 550618 142134 550854
rect 141514 517174 142134 550618
rect 141514 516938 141546 517174
rect 141782 516938 141866 517174
rect 142102 516938 142134 517174
rect 141514 516854 142134 516938
rect 141514 516618 141546 516854
rect 141782 516618 141866 516854
rect 142102 516618 142134 516854
rect 141514 483174 142134 516618
rect 141514 482938 141546 483174
rect 141782 482938 141866 483174
rect 142102 482938 142134 483174
rect 141514 482854 142134 482938
rect 141514 482618 141546 482854
rect 141782 482618 141866 482854
rect 142102 482618 142134 482854
rect 141514 449174 142134 482618
rect 141514 448938 141546 449174
rect 141782 448938 141866 449174
rect 142102 448938 142134 449174
rect 141514 448854 142134 448938
rect 141514 448618 141546 448854
rect 141782 448618 141866 448854
rect 142102 448618 142134 448854
rect 141514 415174 142134 448618
rect 141514 414938 141546 415174
rect 141782 414938 141866 415174
rect 142102 414938 142134 415174
rect 141514 414854 142134 414938
rect 141514 414618 141546 414854
rect 141782 414618 141866 414854
rect 142102 414618 142134 414854
rect 141514 381174 142134 414618
rect 141514 380938 141546 381174
rect 141782 380938 141866 381174
rect 142102 380938 142134 381174
rect 141514 380854 142134 380938
rect 141514 380618 141546 380854
rect 141782 380618 141866 380854
rect 142102 380618 142134 380854
rect 141514 347174 142134 380618
rect 141514 346938 141546 347174
rect 141782 346938 141866 347174
rect 142102 346938 142134 347174
rect 141514 346854 142134 346938
rect 141514 346618 141546 346854
rect 141782 346618 141866 346854
rect 142102 346618 142134 346854
rect 141514 313174 142134 346618
rect 141514 312938 141546 313174
rect 141782 312938 141866 313174
rect 142102 312938 142134 313174
rect 141514 312854 142134 312938
rect 141514 312618 141546 312854
rect 141782 312618 141866 312854
rect 142102 312618 142134 312854
rect 141514 279174 142134 312618
rect 141514 278938 141546 279174
rect 141782 278938 141866 279174
rect 142102 278938 142134 279174
rect 141514 278854 142134 278938
rect 141514 278618 141546 278854
rect 141782 278618 141866 278854
rect 142102 278618 142134 278854
rect 141514 245174 142134 278618
rect 141514 244938 141546 245174
rect 141782 244938 141866 245174
rect 142102 244938 142134 245174
rect 141514 244854 142134 244938
rect 141514 244618 141546 244854
rect 141782 244618 141866 244854
rect 142102 244618 142134 244854
rect 141514 225660 142134 244618
rect 145234 706758 145854 711590
rect 145234 706522 145266 706758
rect 145502 706522 145586 706758
rect 145822 706522 145854 706758
rect 145234 706438 145854 706522
rect 145234 706202 145266 706438
rect 145502 706202 145586 706438
rect 145822 706202 145854 706438
rect 145234 690894 145854 706202
rect 145234 690658 145266 690894
rect 145502 690658 145586 690894
rect 145822 690658 145854 690894
rect 145234 690574 145854 690658
rect 145234 690338 145266 690574
rect 145502 690338 145586 690574
rect 145822 690338 145854 690574
rect 145234 656894 145854 690338
rect 145234 656658 145266 656894
rect 145502 656658 145586 656894
rect 145822 656658 145854 656894
rect 145234 656574 145854 656658
rect 145234 656338 145266 656574
rect 145502 656338 145586 656574
rect 145822 656338 145854 656574
rect 145234 622894 145854 656338
rect 145234 622658 145266 622894
rect 145502 622658 145586 622894
rect 145822 622658 145854 622894
rect 145234 622574 145854 622658
rect 145234 622338 145266 622574
rect 145502 622338 145586 622574
rect 145822 622338 145854 622574
rect 145234 588894 145854 622338
rect 145234 588658 145266 588894
rect 145502 588658 145586 588894
rect 145822 588658 145854 588894
rect 145234 588574 145854 588658
rect 145234 588338 145266 588574
rect 145502 588338 145586 588574
rect 145822 588338 145854 588574
rect 145234 554894 145854 588338
rect 145234 554658 145266 554894
rect 145502 554658 145586 554894
rect 145822 554658 145854 554894
rect 145234 554574 145854 554658
rect 145234 554338 145266 554574
rect 145502 554338 145586 554574
rect 145822 554338 145854 554574
rect 145234 520894 145854 554338
rect 145234 520658 145266 520894
rect 145502 520658 145586 520894
rect 145822 520658 145854 520894
rect 145234 520574 145854 520658
rect 145234 520338 145266 520574
rect 145502 520338 145586 520574
rect 145822 520338 145854 520574
rect 145234 486894 145854 520338
rect 145234 486658 145266 486894
rect 145502 486658 145586 486894
rect 145822 486658 145854 486894
rect 145234 486574 145854 486658
rect 145234 486338 145266 486574
rect 145502 486338 145586 486574
rect 145822 486338 145854 486574
rect 145234 452894 145854 486338
rect 145234 452658 145266 452894
rect 145502 452658 145586 452894
rect 145822 452658 145854 452894
rect 145234 452574 145854 452658
rect 145234 452338 145266 452574
rect 145502 452338 145586 452574
rect 145822 452338 145854 452574
rect 145234 418894 145854 452338
rect 145234 418658 145266 418894
rect 145502 418658 145586 418894
rect 145822 418658 145854 418894
rect 145234 418574 145854 418658
rect 145234 418338 145266 418574
rect 145502 418338 145586 418574
rect 145822 418338 145854 418574
rect 145234 384894 145854 418338
rect 145234 384658 145266 384894
rect 145502 384658 145586 384894
rect 145822 384658 145854 384894
rect 145234 384574 145854 384658
rect 145234 384338 145266 384574
rect 145502 384338 145586 384574
rect 145822 384338 145854 384574
rect 145234 350894 145854 384338
rect 145234 350658 145266 350894
rect 145502 350658 145586 350894
rect 145822 350658 145854 350894
rect 145234 350574 145854 350658
rect 145234 350338 145266 350574
rect 145502 350338 145586 350574
rect 145822 350338 145854 350574
rect 145234 316894 145854 350338
rect 145234 316658 145266 316894
rect 145502 316658 145586 316894
rect 145822 316658 145854 316894
rect 145234 316574 145854 316658
rect 145234 316338 145266 316574
rect 145502 316338 145586 316574
rect 145822 316338 145854 316574
rect 145234 282894 145854 316338
rect 145234 282658 145266 282894
rect 145502 282658 145586 282894
rect 145822 282658 145854 282894
rect 145234 282574 145854 282658
rect 145234 282338 145266 282574
rect 145502 282338 145586 282574
rect 145822 282338 145854 282574
rect 145234 248894 145854 282338
rect 145234 248658 145266 248894
rect 145502 248658 145586 248894
rect 145822 248658 145854 248894
rect 145234 248574 145854 248658
rect 145234 248338 145266 248574
rect 145502 248338 145586 248574
rect 145822 248338 145854 248574
rect 145234 225660 145854 248338
rect 148954 707718 149574 711590
rect 148954 707482 148986 707718
rect 149222 707482 149306 707718
rect 149542 707482 149574 707718
rect 148954 707398 149574 707482
rect 148954 707162 148986 707398
rect 149222 707162 149306 707398
rect 149542 707162 149574 707398
rect 148954 694614 149574 707162
rect 148954 694378 148986 694614
rect 149222 694378 149306 694614
rect 149542 694378 149574 694614
rect 148954 694294 149574 694378
rect 148954 694058 148986 694294
rect 149222 694058 149306 694294
rect 149542 694058 149574 694294
rect 148954 660614 149574 694058
rect 148954 660378 148986 660614
rect 149222 660378 149306 660614
rect 149542 660378 149574 660614
rect 148954 660294 149574 660378
rect 148954 660058 148986 660294
rect 149222 660058 149306 660294
rect 149542 660058 149574 660294
rect 148954 626614 149574 660058
rect 148954 626378 148986 626614
rect 149222 626378 149306 626614
rect 149542 626378 149574 626614
rect 148954 626294 149574 626378
rect 148954 626058 148986 626294
rect 149222 626058 149306 626294
rect 149542 626058 149574 626294
rect 148954 592614 149574 626058
rect 148954 592378 148986 592614
rect 149222 592378 149306 592614
rect 149542 592378 149574 592614
rect 148954 592294 149574 592378
rect 148954 592058 148986 592294
rect 149222 592058 149306 592294
rect 149542 592058 149574 592294
rect 148954 558614 149574 592058
rect 148954 558378 148986 558614
rect 149222 558378 149306 558614
rect 149542 558378 149574 558614
rect 148954 558294 149574 558378
rect 148954 558058 148986 558294
rect 149222 558058 149306 558294
rect 149542 558058 149574 558294
rect 148954 524614 149574 558058
rect 148954 524378 148986 524614
rect 149222 524378 149306 524614
rect 149542 524378 149574 524614
rect 148954 524294 149574 524378
rect 148954 524058 148986 524294
rect 149222 524058 149306 524294
rect 149542 524058 149574 524294
rect 148954 490614 149574 524058
rect 148954 490378 148986 490614
rect 149222 490378 149306 490614
rect 149542 490378 149574 490614
rect 148954 490294 149574 490378
rect 148954 490058 148986 490294
rect 149222 490058 149306 490294
rect 149542 490058 149574 490294
rect 148954 456614 149574 490058
rect 148954 456378 148986 456614
rect 149222 456378 149306 456614
rect 149542 456378 149574 456614
rect 148954 456294 149574 456378
rect 148954 456058 148986 456294
rect 149222 456058 149306 456294
rect 149542 456058 149574 456294
rect 148954 422614 149574 456058
rect 148954 422378 148986 422614
rect 149222 422378 149306 422614
rect 149542 422378 149574 422614
rect 148954 422294 149574 422378
rect 148954 422058 148986 422294
rect 149222 422058 149306 422294
rect 149542 422058 149574 422294
rect 148954 388614 149574 422058
rect 148954 388378 148986 388614
rect 149222 388378 149306 388614
rect 149542 388378 149574 388614
rect 148954 388294 149574 388378
rect 148954 388058 148986 388294
rect 149222 388058 149306 388294
rect 149542 388058 149574 388294
rect 148954 354614 149574 388058
rect 148954 354378 148986 354614
rect 149222 354378 149306 354614
rect 149542 354378 149574 354614
rect 148954 354294 149574 354378
rect 148954 354058 148986 354294
rect 149222 354058 149306 354294
rect 149542 354058 149574 354294
rect 148954 320614 149574 354058
rect 148954 320378 148986 320614
rect 149222 320378 149306 320614
rect 149542 320378 149574 320614
rect 148954 320294 149574 320378
rect 148954 320058 148986 320294
rect 149222 320058 149306 320294
rect 149542 320058 149574 320294
rect 148954 286614 149574 320058
rect 148954 286378 148986 286614
rect 149222 286378 149306 286614
rect 149542 286378 149574 286614
rect 148954 286294 149574 286378
rect 148954 286058 148986 286294
rect 149222 286058 149306 286294
rect 149542 286058 149574 286294
rect 148954 252614 149574 286058
rect 148954 252378 148986 252614
rect 149222 252378 149306 252614
rect 149542 252378 149574 252614
rect 148954 252294 149574 252378
rect 148954 252058 148986 252294
rect 149222 252058 149306 252294
rect 149542 252058 149574 252294
rect 148954 225660 149574 252058
rect 152674 708678 153294 711590
rect 152674 708442 152706 708678
rect 152942 708442 153026 708678
rect 153262 708442 153294 708678
rect 152674 708358 153294 708442
rect 152674 708122 152706 708358
rect 152942 708122 153026 708358
rect 153262 708122 153294 708358
rect 152674 698334 153294 708122
rect 152674 698098 152706 698334
rect 152942 698098 153026 698334
rect 153262 698098 153294 698334
rect 152674 698014 153294 698098
rect 152674 697778 152706 698014
rect 152942 697778 153026 698014
rect 153262 697778 153294 698014
rect 152674 664334 153294 697778
rect 152674 664098 152706 664334
rect 152942 664098 153026 664334
rect 153262 664098 153294 664334
rect 152674 664014 153294 664098
rect 152674 663778 152706 664014
rect 152942 663778 153026 664014
rect 153262 663778 153294 664014
rect 152674 630334 153294 663778
rect 152674 630098 152706 630334
rect 152942 630098 153026 630334
rect 153262 630098 153294 630334
rect 152674 630014 153294 630098
rect 152674 629778 152706 630014
rect 152942 629778 153026 630014
rect 153262 629778 153294 630014
rect 152674 596334 153294 629778
rect 152674 596098 152706 596334
rect 152942 596098 153026 596334
rect 153262 596098 153294 596334
rect 152674 596014 153294 596098
rect 152674 595778 152706 596014
rect 152942 595778 153026 596014
rect 153262 595778 153294 596014
rect 152674 562334 153294 595778
rect 152674 562098 152706 562334
rect 152942 562098 153026 562334
rect 153262 562098 153294 562334
rect 152674 562014 153294 562098
rect 152674 561778 152706 562014
rect 152942 561778 153026 562014
rect 153262 561778 153294 562014
rect 152674 528334 153294 561778
rect 152674 528098 152706 528334
rect 152942 528098 153026 528334
rect 153262 528098 153294 528334
rect 152674 528014 153294 528098
rect 152674 527778 152706 528014
rect 152942 527778 153026 528014
rect 153262 527778 153294 528014
rect 152674 494334 153294 527778
rect 152674 494098 152706 494334
rect 152942 494098 153026 494334
rect 153262 494098 153294 494334
rect 152674 494014 153294 494098
rect 152674 493778 152706 494014
rect 152942 493778 153026 494014
rect 153262 493778 153294 494014
rect 152674 460334 153294 493778
rect 152674 460098 152706 460334
rect 152942 460098 153026 460334
rect 153262 460098 153294 460334
rect 152674 460014 153294 460098
rect 152674 459778 152706 460014
rect 152942 459778 153026 460014
rect 153262 459778 153294 460014
rect 152674 426334 153294 459778
rect 152674 426098 152706 426334
rect 152942 426098 153026 426334
rect 153262 426098 153294 426334
rect 152674 426014 153294 426098
rect 152674 425778 152706 426014
rect 152942 425778 153026 426014
rect 153262 425778 153294 426014
rect 152674 392334 153294 425778
rect 152674 392098 152706 392334
rect 152942 392098 153026 392334
rect 153262 392098 153294 392334
rect 152674 392014 153294 392098
rect 152674 391778 152706 392014
rect 152942 391778 153026 392014
rect 153262 391778 153294 392014
rect 152674 358334 153294 391778
rect 152674 358098 152706 358334
rect 152942 358098 153026 358334
rect 153262 358098 153294 358334
rect 152674 358014 153294 358098
rect 152674 357778 152706 358014
rect 152942 357778 153026 358014
rect 153262 357778 153294 358014
rect 152674 324334 153294 357778
rect 152674 324098 152706 324334
rect 152942 324098 153026 324334
rect 153262 324098 153294 324334
rect 152674 324014 153294 324098
rect 152674 323778 152706 324014
rect 152942 323778 153026 324014
rect 153262 323778 153294 324014
rect 152674 290334 153294 323778
rect 152674 290098 152706 290334
rect 152942 290098 153026 290334
rect 153262 290098 153294 290334
rect 152674 290014 153294 290098
rect 152674 289778 152706 290014
rect 152942 289778 153026 290014
rect 153262 289778 153294 290014
rect 152674 256334 153294 289778
rect 152674 256098 152706 256334
rect 152942 256098 153026 256334
rect 153262 256098 153294 256334
rect 152674 256014 153294 256098
rect 152674 255778 152706 256014
rect 152942 255778 153026 256014
rect 153262 255778 153294 256014
rect 152674 225660 153294 255778
rect 156394 709638 157014 711590
rect 156394 709402 156426 709638
rect 156662 709402 156746 709638
rect 156982 709402 157014 709638
rect 156394 709318 157014 709402
rect 156394 709082 156426 709318
rect 156662 709082 156746 709318
rect 156982 709082 157014 709318
rect 156394 668054 157014 709082
rect 156394 667818 156426 668054
rect 156662 667818 156746 668054
rect 156982 667818 157014 668054
rect 156394 667734 157014 667818
rect 156394 667498 156426 667734
rect 156662 667498 156746 667734
rect 156982 667498 157014 667734
rect 156394 634054 157014 667498
rect 156394 633818 156426 634054
rect 156662 633818 156746 634054
rect 156982 633818 157014 634054
rect 156394 633734 157014 633818
rect 156394 633498 156426 633734
rect 156662 633498 156746 633734
rect 156982 633498 157014 633734
rect 156394 600054 157014 633498
rect 156394 599818 156426 600054
rect 156662 599818 156746 600054
rect 156982 599818 157014 600054
rect 156394 599734 157014 599818
rect 156394 599498 156426 599734
rect 156662 599498 156746 599734
rect 156982 599498 157014 599734
rect 156394 566054 157014 599498
rect 156394 565818 156426 566054
rect 156662 565818 156746 566054
rect 156982 565818 157014 566054
rect 156394 565734 157014 565818
rect 156394 565498 156426 565734
rect 156662 565498 156746 565734
rect 156982 565498 157014 565734
rect 156394 532054 157014 565498
rect 156394 531818 156426 532054
rect 156662 531818 156746 532054
rect 156982 531818 157014 532054
rect 156394 531734 157014 531818
rect 156394 531498 156426 531734
rect 156662 531498 156746 531734
rect 156982 531498 157014 531734
rect 156394 498054 157014 531498
rect 156394 497818 156426 498054
rect 156662 497818 156746 498054
rect 156982 497818 157014 498054
rect 156394 497734 157014 497818
rect 156394 497498 156426 497734
rect 156662 497498 156746 497734
rect 156982 497498 157014 497734
rect 156394 464054 157014 497498
rect 156394 463818 156426 464054
rect 156662 463818 156746 464054
rect 156982 463818 157014 464054
rect 156394 463734 157014 463818
rect 156394 463498 156426 463734
rect 156662 463498 156746 463734
rect 156982 463498 157014 463734
rect 156394 430054 157014 463498
rect 156394 429818 156426 430054
rect 156662 429818 156746 430054
rect 156982 429818 157014 430054
rect 156394 429734 157014 429818
rect 156394 429498 156426 429734
rect 156662 429498 156746 429734
rect 156982 429498 157014 429734
rect 156394 396054 157014 429498
rect 156394 395818 156426 396054
rect 156662 395818 156746 396054
rect 156982 395818 157014 396054
rect 156394 395734 157014 395818
rect 156394 395498 156426 395734
rect 156662 395498 156746 395734
rect 156982 395498 157014 395734
rect 156394 362054 157014 395498
rect 156394 361818 156426 362054
rect 156662 361818 156746 362054
rect 156982 361818 157014 362054
rect 156394 361734 157014 361818
rect 156394 361498 156426 361734
rect 156662 361498 156746 361734
rect 156982 361498 157014 361734
rect 156394 328054 157014 361498
rect 156394 327818 156426 328054
rect 156662 327818 156746 328054
rect 156982 327818 157014 328054
rect 156394 327734 157014 327818
rect 156394 327498 156426 327734
rect 156662 327498 156746 327734
rect 156982 327498 157014 327734
rect 156394 294054 157014 327498
rect 156394 293818 156426 294054
rect 156662 293818 156746 294054
rect 156982 293818 157014 294054
rect 156394 293734 157014 293818
rect 156394 293498 156426 293734
rect 156662 293498 156746 293734
rect 156982 293498 157014 293734
rect 156394 260054 157014 293498
rect 156394 259818 156426 260054
rect 156662 259818 156746 260054
rect 156982 259818 157014 260054
rect 156394 259734 157014 259818
rect 156394 259498 156426 259734
rect 156662 259498 156746 259734
rect 156982 259498 157014 259734
rect 156394 225991 157014 259498
rect 156394 225755 156426 225991
rect 156662 225755 156746 225991
rect 156982 225755 157014 225991
rect 156394 225660 157014 225755
rect 160114 710598 160734 711590
rect 160114 710362 160146 710598
rect 160382 710362 160466 710598
rect 160702 710362 160734 710598
rect 160114 710278 160734 710362
rect 160114 710042 160146 710278
rect 160382 710042 160466 710278
rect 160702 710042 160734 710278
rect 160114 671774 160734 710042
rect 160114 671538 160146 671774
rect 160382 671538 160466 671774
rect 160702 671538 160734 671774
rect 160114 671454 160734 671538
rect 160114 671218 160146 671454
rect 160382 671218 160466 671454
rect 160702 671218 160734 671454
rect 160114 637774 160734 671218
rect 160114 637538 160146 637774
rect 160382 637538 160466 637774
rect 160702 637538 160734 637774
rect 160114 637454 160734 637538
rect 160114 637218 160146 637454
rect 160382 637218 160466 637454
rect 160702 637218 160734 637454
rect 160114 603774 160734 637218
rect 160114 603538 160146 603774
rect 160382 603538 160466 603774
rect 160702 603538 160734 603774
rect 160114 603454 160734 603538
rect 160114 603218 160146 603454
rect 160382 603218 160466 603454
rect 160702 603218 160734 603454
rect 160114 569774 160734 603218
rect 160114 569538 160146 569774
rect 160382 569538 160466 569774
rect 160702 569538 160734 569774
rect 160114 569454 160734 569538
rect 160114 569218 160146 569454
rect 160382 569218 160466 569454
rect 160702 569218 160734 569454
rect 160114 535774 160734 569218
rect 160114 535538 160146 535774
rect 160382 535538 160466 535774
rect 160702 535538 160734 535774
rect 160114 535454 160734 535538
rect 160114 535218 160146 535454
rect 160382 535218 160466 535454
rect 160702 535218 160734 535454
rect 160114 501774 160734 535218
rect 160114 501538 160146 501774
rect 160382 501538 160466 501774
rect 160702 501538 160734 501774
rect 160114 501454 160734 501538
rect 160114 501218 160146 501454
rect 160382 501218 160466 501454
rect 160702 501218 160734 501454
rect 160114 467774 160734 501218
rect 160114 467538 160146 467774
rect 160382 467538 160466 467774
rect 160702 467538 160734 467774
rect 160114 467454 160734 467538
rect 160114 467218 160146 467454
rect 160382 467218 160466 467454
rect 160702 467218 160734 467454
rect 160114 433774 160734 467218
rect 160114 433538 160146 433774
rect 160382 433538 160466 433774
rect 160702 433538 160734 433774
rect 160114 433454 160734 433538
rect 160114 433218 160146 433454
rect 160382 433218 160466 433454
rect 160702 433218 160734 433454
rect 160114 399774 160734 433218
rect 160114 399538 160146 399774
rect 160382 399538 160466 399774
rect 160702 399538 160734 399774
rect 160114 399454 160734 399538
rect 160114 399218 160146 399454
rect 160382 399218 160466 399454
rect 160702 399218 160734 399454
rect 160114 365774 160734 399218
rect 160114 365538 160146 365774
rect 160382 365538 160466 365774
rect 160702 365538 160734 365774
rect 160114 365454 160734 365538
rect 160114 365218 160146 365454
rect 160382 365218 160466 365454
rect 160702 365218 160734 365454
rect 160114 331774 160734 365218
rect 160114 331538 160146 331774
rect 160382 331538 160466 331774
rect 160702 331538 160734 331774
rect 160114 331454 160734 331538
rect 160114 331218 160146 331454
rect 160382 331218 160466 331454
rect 160702 331218 160734 331454
rect 160114 297774 160734 331218
rect 160114 297538 160146 297774
rect 160382 297538 160466 297774
rect 160702 297538 160734 297774
rect 160114 297454 160734 297538
rect 160114 297218 160146 297454
rect 160382 297218 160466 297454
rect 160702 297218 160734 297454
rect 160114 263774 160734 297218
rect 160114 263538 160146 263774
rect 160382 263538 160466 263774
rect 160702 263538 160734 263774
rect 160114 263454 160734 263538
rect 160114 263218 160146 263454
rect 160382 263218 160466 263454
rect 160702 263218 160734 263454
rect 160114 229774 160734 263218
rect 160114 229538 160146 229774
rect 160382 229538 160466 229774
rect 160702 229538 160734 229774
rect 160114 229454 160734 229538
rect 160114 229218 160146 229454
rect 160382 229218 160466 229454
rect 160702 229218 160734 229454
rect 129834 199258 129866 199494
rect 130102 199258 130186 199494
rect 130422 199258 130454 199494
rect 129834 199174 130454 199258
rect 129834 198938 129866 199174
rect 130102 198938 130186 199174
rect 130422 198938 130454 199174
rect 129834 165494 130454 198938
rect 160114 195774 160734 229218
rect 163834 711558 164454 711590
rect 163834 711322 163866 711558
rect 164102 711322 164186 711558
rect 164422 711322 164454 711558
rect 163834 711238 164454 711322
rect 163834 711002 163866 711238
rect 164102 711002 164186 711238
rect 164422 711002 164454 711238
rect 163834 675494 164454 711002
rect 163834 675258 163866 675494
rect 164102 675258 164186 675494
rect 164422 675258 164454 675494
rect 163834 675174 164454 675258
rect 163834 674938 163866 675174
rect 164102 674938 164186 675174
rect 164422 674938 164454 675174
rect 163834 641494 164454 674938
rect 163834 641258 163866 641494
rect 164102 641258 164186 641494
rect 164422 641258 164454 641494
rect 163834 641174 164454 641258
rect 163834 640938 163866 641174
rect 164102 640938 164186 641174
rect 164422 640938 164454 641174
rect 163834 607494 164454 640938
rect 163834 607258 163866 607494
rect 164102 607258 164186 607494
rect 164422 607258 164454 607494
rect 163834 607174 164454 607258
rect 163834 606938 163866 607174
rect 164102 606938 164186 607174
rect 164422 606938 164454 607174
rect 163834 573494 164454 606938
rect 163834 573258 163866 573494
rect 164102 573258 164186 573494
rect 164422 573258 164454 573494
rect 163834 573174 164454 573258
rect 163834 572938 163866 573174
rect 164102 572938 164186 573174
rect 164422 572938 164454 573174
rect 163834 539494 164454 572938
rect 163834 539258 163866 539494
rect 164102 539258 164186 539494
rect 164422 539258 164454 539494
rect 163834 539174 164454 539258
rect 163834 538938 163866 539174
rect 164102 538938 164186 539174
rect 164422 538938 164454 539174
rect 163834 505494 164454 538938
rect 163834 505258 163866 505494
rect 164102 505258 164186 505494
rect 164422 505258 164454 505494
rect 163834 505174 164454 505258
rect 163834 504938 163866 505174
rect 164102 504938 164186 505174
rect 164422 504938 164454 505174
rect 163834 471494 164454 504938
rect 163834 471258 163866 471494
rect 164102 471258 164186 471494
rect 164422 471258 164454 471494
rect 163834 471174 164454 471258
rect 163834 470938 163866 471174
rect 164102 470938 164186 471174
rect 164422 470938 164454 471174
rect 163834 437494 164454 470938
rect 163834 437258 163866 437494
rect 164102 437258 164186 437494
rect 164422 437258 164454 437494
rect 163834 437174 164454 437258
rect 163834 436938 163866 437174
rect 164102 436938 164186 437174
rect 164422 436938 164454 437174
rect 163834 403494 164454 436938
rect 163834 403258 163866 403494
rect 164102 403258 164186 403494
rect 164422 403258 164454 403494
rect 163834 403174 164454 403258
rect 163834 402938 163866 403174
rect 164102 402938 164186 403174
rect 164422 402938 164454 403174
rect 163834 369494 164454 402938
rect 163834 369258 163866 369494
rect 164102 369258 164186 369494
rect 164422 369258 164454 369494
rect 163834 369174 164454 369258
rect 163834 368938 163866 369174
rect 164102 368938 164186 369174
rect 164422 368938 164454 369174
rect 163834 335494 164454 368938
rect 163834 335258 163866 335494
rect 164102 335258 164186 335494
rect 164422 335258 164454 335494
rect 163834 335174 164454 335258
rect 163834 334938 163866 335174
rect 164102 334938 164186 335174
rect 164422 334938 164454 335174
rect 163834 301494 164454 334938
rect 163834 301258 163866 301494
rect 164102 301258 164186 301494
rect 164422 301258 164454 301494
rect 163834 301174 164454 301258
rect 163834 300938 163866 301174
rect 164102 300938 164186 301174
rect 164422 300938 164454 301174
rect 163834 267494 164454 300938
rect 163834 267258 163866 267494
rect 164102 267258 164186 267494
rect 164422 267258 164454 267494
rect 163834 267174 164454 267258
rect 163834 266938 163866 267174
rect 164102 266938 164186 267174
rect 164422 266938 164454 267174
rect 163834 233494 164454 266938
rect 163834 233258 163866 233494
rect 164102 233258 164186 233494
rect 164422 233258 164454 233494
rect 163834 233174 164454 233258
rect 163834 232938 163866 233174
rect 164102 232938 164186 233174
rect 164422 232938 164454 233174
rect 163834 225660 164454 232938
rect 171794 704838 172414 711590
rect 171794 704602 171826 704838
rect 172062 704602 172146 704838
rect 172382 704602 172414 704838
rect 171794 704518 172414 704602
rect 171794 704282 171826 704518
rect 172062 704282 172146 704518
rect 172382 704282 172414 704518
rect 171794 683454 172414 704282
rect 171794 683218 171826 683454
rect 172062 683218 172146 683454
rect 172382 683218 172414 683454
rect 171794 683134 172414 683218
rect 171794 682898 171826 683134
rect 172062 682898 172146 683134
rect 172382 682898 172414 683134
rect 171794 649454 172414 682898
rect 171794 649218 171826 649454
rect 172062 649218 172146 649454
rect 172382 649218 172414 649454
rect 171794 649134 172414 649218
rect 171794 648898 171826 649134
rect 172062 648898 172146 649134
rect 172382 648898 172414 649134
rect 171794 615454 172414 648898
rect 171794 615218 171826 615454
rect 172062 615218 172146 615454
rect 172382 615218 172414 615454
rect 171794 615134 172414 615218
rect 171794 614898 171826 615134
rect 172062 614898 172146 615134
rect 172382 614898 172414 615134
rect 171794 581454 172414 614898
rect 171794 581218 171826 581454
rect 172062 581218 172146 581454
rect 172382 581218 172414 581454
rect 171794 581134 172414 581218
rect 171794 580898 171826 581134
rect 172062 580898 172146 581134
rect 172382 580898 172414 581134
rect 171794 547454 172414 580898
rect 171794 547218 171826 547454
rect 172062 547218 172146 547454
rect 172382 547218 172414 547454
rect 171794 547134 172414 547218
rect 171794 546898 171826 547134
rect 172062 546898 172146 547134
rect 172382 546898 172414 547134
rect 171794 513454 172414 546898
rect 171794 513218 171826 513454
rect 172062 513218 172146 513454
rect 172382 513218 172414 513454
rect 171794 513134 172414 513218
rect 171794 512898 171826 513134
rect 172062 512898 172146 513134
rect 172382 512898 172414 513134
rect 171794 479454 172414 512898
rect 171794 479218 171826 479454
rect 172062 479218 172146 479454
rect 172382 479218 172414 479454
rect 171794 479134 172414 479218
rect 171794 478898 171826 479134
rect 172062 478898 172146 479134
rect 172382 478898 172414 479134
rect 171794 445454 172414 478898
rect 171794 445218 171826 445454
rect 172062 445218 172146 445454
rect 172382 445218 172414 445454
rect 171794 445134 172414 445218
rect 171794 444898 171826 445134
rect 172062 444898 172146 445134
rect 172382 444898 172414 445134
rect 171794 411454 172414 444898
rect 171794 411218 171826 411454
rect 172062 411218 172146 411454
rect 172382 411218 172414 411454
rect 171794 411134 172414 411218
rect 171794 410898 171826 411134
rect 172062 410898 172146 411134
rect 172382 410898 172414 411134
rect 171794 377454 172414 410898
rect 171794 377218 171826 377454
rect 172062 377218 172146 377454
rect 172382 377218 172414 377454
rect 171794 377134 172414 377218
rect 171794 376898 171826 377134
rect 172062 376898 172146 377134
rect 172382 376898 172414 377134
rect 171794 343454 172414 376898
rect 171794 343218 171826 343454
rect 172062 343218 172146 343454
rect 172382 343218 172414 343454
rect 171794 343134 172414 343218
rect 171794 342898 171826 343134
rect 172062 342898 172146 343134
rect 172382 342898 172414 343134
rect 171794 309454 172414 342898
rect 171794 309218 171826 309454
rect 172062 309218 172146 309454
rect 172382 309218 172414 309454
rect 171794 309134 172414 309218
rect 171794 308898 171826 309134
rect 172062 308898 172146 309134
rect 172382 308898 172414 309134
rect 171794 275454 172414 308898
rect 171794 275218 171826 275454
rect 172062 275218 172146 275454
rect 172382 275218 172414 275454
rect 171794 275134 172414 275218
rect 171794 274898 171826 275134
rect 172062 274898 172146 275134
rect 172382 274898 172414 275134
rect 171794 241454 172414 274898
rect 171794 241218 171826 241454
rect 172062 241218 172146 241454
rect 172382 241218 172414 241454
rect 171794 241134 172414 241218
rect 171794 240898 171826 241134
rect 172062 240898 172146 241134
rect 172382 240898 172414 241134
rect 171794 225660 172414 240898
rect 175514 705798 176134 711590
rect 175514 705562 175546 705798
rect 175782 705562 175866 705798
rect 176102 705562 176134 705798
rect 175514 705478 176134 705562
rect 175514 705242 175546 705478
rect 175782 705242 175866 705478
rect 176102 705242 176134 705478
rect 175514 687174 176134 705242
rect 175514 686938 175546 687174
rect 175782 686938 175866 687174
rect 176102 686938 176134 687174
rect 175514 686854 176134 686938
rect 175514 686618 175546 686854
rect 175782 686618 175866 686854
rect 176102 686618 176134 686854
rect 175514 653174 176134 686618
rect 175514 652938 175546 653174
rect 175782 652938 175866 653174
rect 176102 652938 176134 653174
rect 175514 652854 176134 652938
rect 175514 652618 175546 652854
rect 175782 652618 175866 652854
rect 176102 652618 176134 652854
rect 175514 619174 176134 652618
rect 175514 618938 175546 619174
rect 175782 618938 175866 619174
rect 176102 618938 176134 619174
rect 175514 618854 176134 618938
rect 175514 618618 175546 618854
rect 175782 618618 175866 618854
rect 176102 618618 176134 618854
rect 175514 585174 176134 618618
rect 175514 584938 175546 585174
rect 175782 584938 175866 585174
rect 176102 584938 176134 585174
rect 175514 584854 176134 584938
rect 175514 584618 175546 584854
rect 175782 584618 175866 584854
rect 176102 584618 176134 584854
rect 175514 551174 176134 584618
rect 175514 550938 175546 551174
rect 175782 550938 175866 551174
rect 176102 550938 176134 551174
rect 175514 550854 176134 550938
rect 175514 550618 175546 550854
rect 175782 550618 175866 550854
rect 176102 550618 176134 550854
rect 175514 517174 176134 550618
rect 175514 516938 175546 517174
rect 175782 516938 175866 517174
rect 176102 516938 176134 517174
rect 175514 516854 176134 516938
rect 175514 516618 175546 516854
rect 175782 516618 175866 516854
rect 176102 516618 176134 516854
rect 175514 483174 176134 516618
rect 175514 482938 175546 483174
rect 175782 482938 175866 483174
rect 176102 482938 176134 483174
rect 175514 482854 176134 482938
rect 175514 482618 175546 482854
rect 175782 482618 175866 482854
rect 176102 482618 176134 482854
rect 175514 449174 176134 482618
rect 175514 448938 175546 449174
rect 175782 448938 175866 449174
rect 176102 448938 176134 449174
rect 175514 448854 176134 448938
rect 175514 448618 175546 448854
rect 175782 448618 175866 448854
rect 176102 448618 176134 448854
rect 175514 415174 176134 448618
rect 175514 414938 175546 415174
rect 175782 414938 175866 415174
rect 176102 414938 176134 415174
rect 175514 414854 176134 414938
rect 175514 414618 175546 414854
rect 175782 414618 175866 414854
rect 176102 414618 176134 414854
rect 175514 381174 176134 414618
rect 175514 380938 175546 381174
rect 175782 380938 175866 381174
rect 176102 380938 176134 381174
rect 175514 380854 176134 380938
rect 175514 380618 175546 380854
rect 175782 380618 175866 380854
rect 176102 380618 176134 380854
rect 175514 347174 176134 380618
rect 175514 346938 175546 347174
rect 175782 346938 175866 347174
rect 176102 346938 176134 347174
rect 175514 346854 176134 346938
rect 175514 346618 175546 346854
rect 175782 346618 175866 346854
rect 176102 346618 176134 346854
rect 175514 313174 176134 346618
rect 175514 312938 175546 313174
rect 175782 312938 175866 313174
rect 176102 312938 176134 313174
rect 175514 312854 176134 312938
rect 175514 312618 175546 312854
rect 175782 312618 175866 312854
rect 176102 312618 176134 312854
rect 175514 279174 176134 312618
rect 175514 278938 175546 279174
rect 175782 278938 175866 279174
rect 176102 278938 176134 279174
rect 175514 278854 176134 278938
rect 175514 278618 175546 278854
rect 175782 278618 175866 278854
rect 176102 278618 176134 278854
rect 175514 245174 176134 278618
rect 175514 244938 175546 245174
rect 175782 244938 175866 245174
rect 176102 244938 176134 245174
rect 175514 244854 176134 244938
rect 175514 244618 175546 244854
rect 175782 244618 175866 244854
rect 176102 244618 176134 244854
rect 175514 225660 176134 244618
rect 179234 706758 179854 711590
rect 179234 706522 179266 706758
rect 179502 706522 179586 706758
rect 179822 706522 179854 706758
rect 179234 706438 179854 706522
rect 179234 706202 179266 706438
rect 179502 706202 179586 706438
rect 179822 706202 179854 706438
rect 179234 690894 179854 706202
rect 179234 690658 179266 690894
rect 179502 690658 179586 690894
rect 179822 690658 179854 690894
rect 179234 690574 179854 690658
rect 179234 690338 179266 690574
rect 179502 690338 179586 690574
rect 179822 690338 179854 690574
rect 179234 656894 179854 690338
rect 179234 656658 179266 656894
rect 179502 656658 179586 656894
rect 179822 656658 179854 656894
rect 179234 656574 179854 656658
rect 179234 656338 179266 656574
rect 179502 656338 179586 656574
rect 179822 656338 179854 656574
rect 179234 622894 179854 656338
rect 179234 622658 179266 622894
rect 179502 622658 179586 622894
rect 179822 622658 179854 622894
rect 179234 622574 179854 622658
rect 179234 622338 179266 622574
rect 179502 622338 179586 622574
rect 179822 622338 179854 622574
rect 179234 588894 179854 622338
rect 179234 588658 179266 588894
rect 179502 588658 179586 588894
rect 179822 588658 179854 588894
rect 179234 588574 179854 588658
rect 179234 588338 179266 588574
rect 179502 588338 179586 588574
rect 179822 588338 179854 588574
rect 179234 554894 179854 588338
rect 179234 554658 179266 554894
rect 179502 554658 179586 554894
rect 179822 554658 179854 554894
rect 179234 554574 179854 554658
rect 179234 554338 179266 554574
rect 179502 554338 179586 554574
rect 179822 554338 179854 554574
rect 179234 520894 179854 554338
rect 179234 520658 179266 520894
rect 179502 520658 179586 520894
rect 179822 520658 179854 520894
rect 179234 520574 179854 520658
rect 179234 520338 179266 520574
rect 179502 520338 179586 520574
rect 179822 520338 179854 520574
rect 179234 486894 179854 520338
rect 179234 486658 179266 486894
rect 179502 486658 179586 486894
rect 179822 486658 179854 486894
rect 179234 486574 179854 486658
rect 179234 486338 179266 486574
rect 179502 486338 179586 486574
rect 179822 486338 179854 486574
rect 179234 452894 179854 486338
rect 179234 452658 179266 452894
rect 179502 452658 179586 452894
rect 179822 452658 179854 452894
rect 179234 452574 179854 452658
rect 179234 452338 179266 452574
rect 179502 452338 179586 452574
rect 179822 452338 179854 452574
rect 179234 418894 179854 452338
rect 179234 418658 179266 418894
rect 179502 418658 179586 418894
rect 179822 418658 179854 418894
rect 179234 418574 179854 418658
rect 179234 418338 179266 418574
rect 179502 418338 179586 418574
rect 179822 418338 179854 418574
rect 179234 384894 179854 418338
rect 179234 384658 179266 384894
rect 179502 384658 179586 384894
rect 179822 384658 179854 384894
rect 179234 384574 179854 384658
rect 179234 384338 179266 384574
rect 179502 384338 179586 384574
rect 179822 384338 179854 384574
rect 179234 350894 179854 384338
rect 179234 350658 179266 350894
rect 179502 350658 179586 350894
rect 179822 350658 179854 350894
rect 179234 350574 179854 350658
rect 179234 350338 179266 350574
rect 179502 350338 179586 350574
rect 179822 350338 179854 350574
rect 179234 316894 179854 350338
rect 179234 316658 179266 316894
rect 179502 316658 179586 316894
rect 179822 316658 179854 316894
rect 179234 316574 179854 316658
rect 179234 316338 179266 316574
rect 179502 316338 179586 316574
rect 179822 316338 179854 316574
rect 179234 282894 179854 316338
rect 179234 282658 179266 282894
rect 179502 282658 179586 282894
rect 179822 282658 179854 282894
rect 179234 282574 179854 282658
rect 179234 282338 179266 282574
rect 179502 282338 179586 282574
rect 179822 282338 179854 282574
rect 179234 248894 179854 282338
rect 179234 248658 179266 248894
rect 179502 248658 179586 248894
rect 179822 248658 179854 248894
rect 179234 248574 179854 248658
rect 179234 248338 179266 248574
rect 179502 248338 179586 248574
rect 179822 248338 179854 248574
rect 179234 225660 179854 248338
rect 182954 707718 183574 711590
rect 182954 707482 182986 707718
rect 183222 707482 183306 707718
rect 183542 707482 183574 707718
rect 182954 707398 183574 707482
rect 182954 707162 182986 707398
rect 183222 707162 183306 707398
rect 183542 707162 183574 707398
rect 182954 694614 183574 707162
rect 182954 694378 182986 694614
rect 183222 694378 183306 694614
rect 183542 694378 183574 694614
rect 182954 694294 183574 694378
rect 182954 694058 182986 694294
rect 183222 694058 183306 694294
rect 183542 694058 183574 694294
rect 182954 660614 183574 694058
rect 182954 660378 182986 660614
rect 183222 660378 183306 660614
rect 183542 660378 183574 660614
rect 182954 660294 183574 660378
rect 182954 660058 182986 660294
rect 183222 660058 183306 660294
rect 183542 660058 183574 660294
rect 182954 626614 183574 660058
rect 182954 626378 182986 626614
rect 183222 626378 183306 626614
rect 183542 626378 183574 626614
rect 182954 626294 183574 626378
rect 182954 626058 182986 626294
rect 183222 626058 183306 626294
rect 183542 626058 183574 626294
rect 182954 592614 183574 626058
rect 182954 592378 182986 592614
rect 183222 592378 183306 592614
rect 183542 592378 183574 592614
rect 182954 592294 183574 592378
rect 182954 592058 182986 592294
rect 183222 592058 183306 592294
rect 183542 592058 183574 592294
rect 182954 558614 183574 592058
rect 182954 558378 182986 558614
rect 183222 558378 183306 558614
rect 183542 558378 183574 558614
rect 182954 558294 183574 558378
rect 182954 558058 182986 558294
rect 183222 558058 183306 558294
rect 183542 558058 183574 558294
rect 182954 524614 183574 558058
rect 182954 524378 182986 524614
rect 183222 524378 183306 524614
rect 183542 524378 183574 524614
rect 182954 524294 183574 524378
rect 182954 524058 182986 524294
rect 183222 524058 183306 524294
rect 183542 524058 183574 524294
rect 182954 490614 183574 524058
rect 182954 490378 182986 490614
rect 183222 490378 183306 490614
rect 183542 490378 183574 490614
rect 182954 490294 183574 490378
rect 182954 490058 182986 490294
rect 183222 490058 183306 490294
rect 183542 490058 183574 490294
rect 182954 456614 183574 490058
rect 182954 456378 182986 456614
rect 183222 456378 183306 456614
rect 183542 456378 183574 456614
rect 182954 456294 183574 456378
rect 182954 456058 182986 456294
rect 183222 456058 183306 456294
rect 183542 456058 183574 456294
rect 182954 422614 183574 456058
rect 182954 422378 182986 422614
rect 183222 422378 183306 422614
rect 183542 422378 183574 422614
rect 182954 422294 183574 422378
rect 182954 422058 182986 422294
rect 183222 422058 183306 422294
rect 183542 422058 183574 422294
rect 182954 388614 183574 422058
rect 182954 388378 182986 388614
rect 183222 388378 183306 388614
rect 183542 388378 183574 388614
rect 182954 388294 183574 388378
rect 182954 388058 182986 388294
rect 183222 388058 183306 388294
rect 183542 388058 183574 388294
rect 182954 354614 183574 388058
rect 182954 354378 182986 354614
rect 183222 354378 183306 354614
rect 183542 354378 183574 354614
rect 182954 354294 183574 354378
rect 182954 354058 182986 354294
rect 183222 354058 183306 354294
rect 183542 354058 183574 354294
rect 182954 320614 183574 354058
rect 182954 320378 182986 320614
rect 183222 320378 183306 320614
rect 183542 320378 183574 320614
rect 182954 320294 183574 320378
rect 182954 320058 182986 320294
rect 183222 320058 183306 320294
rect 183542 320058 183574 320294
rect 182954 286614 183574 320058
rect 182954 286378 182986 286614
rect 183222 286378 183306 286614
rect 183542 286378 183574 286614
rect 182954 286294 183574 286378
rect 182954 286058 182986 286294
rect 183222 286058 183306 286294
rect 183542 286058 183574 286294
rect 182954 252614 183574 286058
rect 182954 252378 182986 252614
rect 183222 252378 183306 252614
rect 183542 252378 183574 252614
rect 182954 252294 183574 252378
rect 182954 252058 182986 252294
rect 183222 252058 183306 252294
rect 183542 252058 183574 252294
rect 182954 225660 183574 252058
rect 186674 708678 187294 711590
rect 186674 708442 186706 708678
rect 186942 708442 187026 708678
rect 187262 708442 187294 708678
rect 186674 708358 187294 708442
rect 186674 708122 186706 708358
rect 186942 708122 187026 708358
rect 187262 708122 187294 708358
rect 186674 698334 187294 708122
rect 186674 698098 186706 698334
rect 186942 698098 187026 698334
rect 187262 698098 187294 698334
rect 186674 698014 187294 698098
rect 186674 697778 186706 698014
rect 186942 697778 187026 698014
rect 187262 697778 187294 698014
rect 186674 664334 187294 697778
rect 186674 664098 186706 664334
rect 186942 664098 187026 664334
rect 187262 664098 187294 664334
rect 186674 664014 187294 664098
rect 186674 663778 186706 664014
rect 186942 663778 187026 664014
rect 187262 663778 187294 664014
rect 186674 630334 187294 663778
rect 186674 630098 186706 630334
rect 186942 630098 187026 630334
rect 187262 630098 187294 630334
rect 186674 630014 187294 630098
rect 186674 629778 186706 630014
rect 186942 629778 187026 630014
rect 187262 629778 187294 630014
rect 186674 596334 187294 629778
rect 186674 596098 186706 596334
rect 186942 596098 187026 596334
rect 187262 596098 187294 596334
rect 186674 596014 187294 596098
rect 186674 595778 186706 596014
rect 186942 595778 187026 596014
rect 187262 595778 187294 596014
rect 186674 562334 187294 595778
rect 186674 562098 186706 562334
rect 186942 562098 187026 562334
rect 187262 562098 187294 562334
rect 186674 562014 187294 562098
rect 186674 561778 186706 562014
rect 186942 561778 187026 562014
rect 187262 561778 187294 562014
rect 186674 528334 187294 561778
rect 186674 528098 186706 528334
rect 186942 528098 187026 528334
rect 187262 528098 187294 528334
rect 186674 528014 187294 528098
rect 186674 527778 186706 528014
rect 186942 527778 187026 528014
rect 187262 527778 187294 528014
rect 186674 494334 187294 527778
rect 186674 494098 186706 494334
rect 186942 494098 187026 494334
rect 187262 494098 187294 494334
rect 186674 494014 187294 494098
rect 186674 493778 186706 494014
rect 186942 493778 187026 494014
rect 187262 493778 187294 494014
rect 186674 460334 187294 493778
rect 186674 460098 186706 460334
rect 186942 460098 187026 460334
rect 187262 460098 187294 460334
rect 186674 460014 187294 460098
rect 186674 459778 186706 460014
rect 186942 459778 187026 460014
rect 187262 459778 187294 460014
rect 186674 426334 187294 459778
rect 186674 426098 186706 426334
rect 186942 426098 187026 426334
rect 187262 426098 187294 426334
rect 186674 426014 187294 426098
rect 186674 425778 186706 426014
rect 186942 425778 187026 426014
rect 187262 425778 187294 426014
rect 186674 392334 187294 425778
rect 186674 392098 186706 392334
rect 186942 392098 187026 392334
rect 187262 392098 187294 392334
rect 186674 392014 187294 392098
rect 186674 391778 186706 392014
rect 186942 391778 187026 392014
rect 187262 391778 187294 392014
rect 186674 358334 187294 391778
rect 186674 358098 186706 358334
rect 186942 358098 187026 358334
rect 187262 358098 187294 358334
rect 186674 358014 187294 358098
rect 186674 357778 186706 358014
rect 186942 357778 187026 358014
rect 187262 357778 187294 358014
rect 186674 324334 187294 357778
rect 186674 324098 186706 324334
rect 186942 324098 187026 324334
rect 187262 324098 187294 324334
rect 186674 324014 187294 324098
rect 186674 323778 186706 324014
rect 186942 323778 187026 324014
rect 187262 323778 187294 324014
rect 186674 290334 187294 323778
rect 186674 290098 186706 290334
rect 186942 290098 187026 290334
rect 187262 290098 187294 290334
rect 186674 290014 187294 290098
rect 186674 289778 186706 290014
rect 186942 289778 187026 290014
rect 187262 289778 187294 290014
rect 186674 256334 187294 289778
rect 186674 256098 186706 256334
rect 186942 256098 187026 256334
rect 187262 256098 187294 256334
rect 186674 256014 187294 256098
rect 186674 255778 186706 256014
rect 186942 255778 187026 256014
rect 187262 255778 187294 256014
rect 186674 225660 187294 255778
rect 190394 709638 191014 711590
rect 190394 709402 190426 709638
rect 190662 709402 190746 709638
rect 190982 709402 191014 709638
rect 190394 709318 191014 709402
rect 190394 709082 190426 709318
rect 190662 709082 190746 709318
rect 190982 709082 191014 709318
rect 190394 668054 191014 709082
rect 190394 667818 190426 668054
rect 190662 667818 190746 668054
rect 190982 667818 191014 668054
rect 190394 667734 191014 667818
rect 190394 667498 190426 667734
rect 190662 667498 190746 667734
rect 190982 667498 191014 667734
rect 190394 634054 191014 667498
rect 190394 633818 190426 634054
rect 190662 633818 190746 634054
rect 190982 633818 191014 634054
rect 190394 633734 191014 633818
rect 190394 633498 190426 633734
rect 190662 633498 190746 633734
rect 190982 633498 191014 633734
rect 190394 600054 191014 633498
rect 190394 599818 190426 600054
rect 190662 599818 190746 600054
rect 190982 599818 191014 600054
rect 190394 599734 191014 599818
rect 190394 599498 190426 599734
rect 190662 599498 190746 599734
rect 190982 599498 191014 599734
rect 190394 566054 191014 599498
rect 190394 565818 190426 566054
rect 190662 565818 190746 566054
rect 190982 565818 191014 566054
rect 190394 565734 191014 565818
rect 190394 565498 190426 565734
rect 190662 565498 190746 565734
rect 190982 565498 191014 565734
rect 190394 532054 191014 565498
rect 190394 531818 190426 532054
rect 190662 531818 190746 532054
rect 190982 531818 191014 532054
rect 190394 531734 191014 531818
rect 190394 531498 190426 531734
rect 190662 531498 190746 531734
rect 190982 531498 191014 531734
rect 190394 498054 191014 531498
rect 190394 497818 190426 498054
rect 190662 497818 190746 498054
rect 190982 497818 191014 498054
rect 190394 497734 191014 497818
rect 190394 497498 190426 497734
rect 190662 497498 190746 497734
rect 190982 497498 191014 497734
rect 190394 464054 191014 497498
rect 190394 463818 190426 464054
rect 190662 463818 190746 464054
rect 190982 463818 191014 464054
rect 190394 463734 191014 463818
rect 190394 463498 190426 463734
rect 190662 463498 190746 463734
rect 190982 463498 191014 463734
rect 190394 430054 191014 463498
rect 190394 429818 190426 430054
rect 190662 429818 190746 430054
rect 190982 429818 191014 430054
rect 190394 429734 191014 429818
rect 190394 429498 190426 429734
rect 190662 429498 190746 429734
rect 190982 429498 191014 429734
rect 190394 396054 191014 429498
rect 190394 395818 190426 396054
rect 190662 395818 190746 396054
rect 190982 395818 191014 396054
rect 190394 395734 191014 395818
rect 190394 395498 190426 395734
rect 190662 395498 190746 395734
rect 190982 395498 191014 395734
rect 190394 362054 191014 395498
rect 190394 361818 190426 362054
rect 190662 361818 190746 362054
rect 190982 361818 191014 362054
rect 190394 361734 191014 361818
rect 190394 361498 190426 361734
rect 190662 361498 190746 361734
rect 190982 361498 191014 361734
rect 190394 328054 191014 361498
rect 190394 327818 190426 328054
rect 190662 327818 190746 328054
rect 190982 327818 191014 328054
rect 190394 327734 191014 327818
rect 190394 327498 190426 327734
rect 190662 327498 190746 327734
rect 190982 327498 191014 327734
rect 190394 294054 191014 327498
rect 190394 293818 190426 294054
rect 190662 293818 190746 294054
rect 190982 293818 191014 294054
rect 190394 293734 191014 293818
rect 190394 293498 190426 293734
rect 190662 293498 190746 293734
rect 190982 293498 191014 293734
rect 190394 260054 191014 293498
rect 190394 259818 190426 260054
rect 190662 259818 190746 260054
rect 190982 259818 191014 260054
rect 190394 259734 191014 259818
rect 190394 259498 190426 259734
rect 190662 259498 190746 259734
rect 190982 259498 191014 259734
rect 190394 226054 191014 259498
rect 190394 225818 190426 226054
rect 190662 225818 190746 226054
rect 190982 225818 191014 226054
rect 190394 225734 191014 225818
rect 190394 225498 190426 225734
rect 190662 225498 190746 225734
rect 190982 225498 191014 225734
rect 194114 710598 194734 711590
rect 194114 710362 194146 710598
rect 194382 710362 194466 710598
rect 194702 710362 194734 710598
rect 194114 710278 194734 710362
rect 194114 710042 194146 710278
rect 194382 710042 194466 710278
rect 194702 710042 194734 710278
rect 194114 671774 194734 710042
rect 194114 671538 194146 671774
rect 194382 671538 194466 671774
rect 194702 671538 194734 671774
rect 194114 671454 194734 671538
rect 194114 671218 194146 671454
rect 194382 671218 194466 671454
rect 194702 671218 194734 671454
rect 194114 637774 194734 671218
rect 194114 637538 194146 637774
rect 194382 637538 194466 637774
rect 194702 637538 194734 637774
rect 194114 637454 194734 637538
rect 194114 637218 194146 637454
rect 194382 637218 194466 637454
rect 194702 637218 194734 637454
rect 194114 603774 194734 637218
rect 194114 603538 194146 603774
rect 194382 603538 194466 603774
rect 194702 603538 194734 603774
rect 194114 603454 194734 603538
rect 194114 603218 194146 603454
rect 194382 603218 194466 603454
rect 194702 603218 194734 603454
rect 194114 569774 194734 603218
rect 194114 569538 194146 569774
rect 194382 569538 194466 569774
rect 194702 569538 194734 569774
rect 194114 569454 194734 569538
rect 194114 569218 194146 569454
rect 194382 569218 194466 569454
rect 194702 569218 194734 569454
rect 194114 535774 194734 569218
rect 194114 535538 194146 535774
rect 194382 535538 194466 535774
rect 194702 535538 194734 535774
rect 194114 535454 194734 535538
rect 194114 535218 194146 535454
rect 194382 535218 194466 535454
rect 194702 535218 194734 535454
rect 194114 501774 194734 535218
rect 194114 501538 194146 501774
rect 194382 501538 194466 501774
rect 194702 501538 194734 501774
rect 194114 501454 194734 501538
rect 194114 501218 194146 501454
rect 194382 501218 194466 501454
rect 194702 501218 194734 501454
rect 194114 467774 194734 501218
rect 194114 467538 194146 467774
rect 194382 467538 194466 467774
rect 194702 467538 194734 467774
rect 194114 467454 194734 467538
rect 194114 467218 194146 467454
rect 194382 467218 194466 467454
rect 194702 467218 194734 467454
rect 194114 433774 194734 467218
rect 194114 433538 194146 433774
rect 194382 433538 194466 433774
rect 194702 433538 194734 433774
rect 194114 433454 194734 433538
rect 194114 433218 194146 433454
rect 194382 433218 194466 433454
rect 194702 433218 194734 433454
rect 194114 399774 194734 433218
rect 194114 399538 194146 399774
rect 194382 399538 194466 399774
rect 194702 399538 194734 399774
rect 194114 399454 194734 399538
rect 194114 399218 194146 399454
rect 194382 399218 194466 399454
rect 194702 399218 194734 399454
rect 194114 365774 194734 399218
rect 194114 365538 194146 365774
rect 194382 365538 194466 365774
rect 194702 365538 194734 365774
rect 194114 365454 194734 365538
rect 194114 365218 194146 365454
rect 194382 365218 194466 365454
rect 194702 365218 194734 365454
rect 194114 331774 194734 365218
rect 194114 331538 194146 331774
rect 194382 331538 194466 331774
rect 194702 331538 194734 331774
rect 194114 331454 194734 331538
rect 194114 331218 194146 331454
rect 194382 331218 194466 331454
rect 194702 331218 194734 331454
rect 194114 297774 194734 331218
rect 194114 297538 194146 297774
rect 194382 297538 194466 297774
rect 194702 297538 194734 297774
rect 194114 297454 194734 297538
rect 194114 297218 194146 297454
rect 194382 297218 194466 297454
rect 194702 297218 194734 297454
rect 194114 263774 194734 297218
rect 194114 263538 194146 263774
rect 194382 263538 194466 263774
rect 194702 263538 194734 263774
rect 194114 263454 194734 263538
rect 194114 263218 194146 263454
rect 194382 263218 194466 263454
rect 194702 263218 194734 263454
rect 194114 229774 194734 263218
rect 194114 229538 194146 229774
rect 194382 229538 194466 229774
rect 194702 229538 194734 229774
rect 194114 229454 194734 229538
rect 194114 229218 194146 229454
rect 194382 229218 194466 229454
rect 194702 229218 194734 229454
rect 194114 225660 194734 229218
rect 197834 711558 198454 711590
rect 197834 711322 197866 711558
rect 198102 711322 198186 711558
rect 198422 711322 198454 711558
rect 197834 711238 198454 711322
rect 197834 711002 197866 711238
rect 198102 711002 198186 711238
rect 198422 711002 198454 711238
rect 197834 675494 198454 711002
rect 197834 675258 197866 675494
rect 198102 675258 198186 675494
rect 198422 675258 198454 675494
rect 197834 675174 198454 675258
rect 197834 674938 197866 675174
rect 198102 674938 198186 675174
rect 198422 674938 198454 675174
rect 197834 641494 198454 674938
rect 197834 641258 197866 641494
rect 198102 641258 198186 641494
rect 198422 641258 198454 641494
rect 197834 641174 198454 641258
rect 197834 640938 197866 641174
rect 198102 640938 198186 641174
rect 198422 640938 198454 641174
rect 197834 607494 198454 640938
rect 197834 607258 197866 607494
rect 198102 607258 198186 607494
rect 198422 607258 198454 607494
rect 197834 607174 198454 607258
rect 197834 606938 197866 607174
rect 198102 606938 198186 607174
rect 198422 606938 198454 607174
rect 197834 573494 198454 606938
rect 197834 573258 197866 573494
rect 198102 573258 198186 573494
rect 198422 573258 198454 573494
rect 197834 573174 198454 573258
rect 197834 572938 197866 573174
rect 198102 572938 198186 573174
rect 198422 572938 198454 573174
rect 197834 539494 198454 572938
rect 197834 539258 197866 539494
rect 198102 539258 198186 539494
rect 198422 539258 198454 539494
rect 197834 539174 198454 539258
rect 197834 538938 197866 539174
rect 198102 538938 198186 539174
rect 198422 538938 198454 539174
rect 197834 505494 198454 538938
rect 197834 505258 197866 505494
rect 198102 505258 198186 505494
rect 198422 505258 198454 505494
rect 197834 505174 198454 505258
rect 197834 504938 197866 505174
rect 198102 504938 198186 505174
rect 198422 504938 198454 505174
rect 197834 471494 198454 504938
rect 197834 471258 197866 471494
rect 198102 471258 198186 471494
rect 198422 471258 198454 471494
rect 197834 471174 198454 471258
rect 197834 470938 197866 471174
rect 198102 470938 198186 471174
rect 198422 470938 198454 471174
rect 197834 437494 198454 470938
rect 197834 437258 197866 437494
rect 198102 437258 198186 437494
rect 198422 437258 198454 437494
rect 197834 437174 198454 437258
rect 197834 436938 197866 437174
rect 198102 436938 198186 437174
rect 198422 436938 198454 437174
rect 197834 403494 198454 436938
rect 197834 403258 197866 403494
rect 198102 403258 198186 403494
rect 198422 403258 198454 403494
rect 197834 403174 198454 403258
rect 197834 402938 197866 403174
rect 198102 402938 198186 403174
rect 198422 402938 198454 403174
rect 197834 369494 198454 402938
rect 197834 369258 197866 369494
rect 198102 369258 198186 369494
rect 198422 369258 198454 369494
rect 197834 369174 198454 369258
rect 197834 368938 197866 369174
rect 198102 368938 198186 369174
rect 198422 368938 198454 369174
rect 197834 335494 198454 368938
rect 197834 335258 197866 335494
rect 198102 335258 198186 335494
rect 198422 335258 198454 335494
rect 197834 335174 198454 335258
rect 197834 334938 197866 335174
rect 198102 334938 198186 335174
rect 198422 334938 198454 335174
rect 197834 301494 198454 334938
rect 197834 301258 197866 301494
rect 198102 301258 198186 301494
rect 198422 301258 198454 301494
rect 197834 301174 198454 301258
rect 197834 300938 197866 301174
rect 198102 300938 198186 301174
rect 198422 300938 198454 301174
rect 197834 267494 198454 300938
rect 197834 267258 197866 267494
rect 198102 267258 198186 267494
rect 198422 267258 198454 267494
rect 197834 267174 198454 267258
rect 197834 266938 197866 267174
rect 198102 266938 198186 267174
rect 198422 266938 198454 267174
rect 197834 233494 198454 266938
rect 197834 233258 197866 233494
rect 198102 233258 198186 233494
rect 198422 233258 198454 233494
rect 197834 233174 198454 233258
rect 197834 232938 197866 233174
rect 198102 232938 198186 233174
rect 198422 232938 198454 233174
rect 197834 225660 198454 232938
rect 205794 704838 206414 711590
rect 205794 704602 205826 704838
rect 206062 704602 206146 704838
rect 206382 704602 206414 704838
rect 205794 704518 206414 704602
rect 205794 704282 205826 704518
rect 206062 704282 206146 704518
rect 206382 704282 206414 704518
rect 205794 683454 206414 704282
rect 205794 683218 205826 683454
rect 206062 683218 206146 683454
rect 206382 683218 206414 683454
rect 205794 683134 206414 683218
rect 205794 682898 205826 683134
rect 206062 682898 206146 683134
rect 206382 682898 206414 683134
rect 205794 649454 206414 682898
rect 205794 649218 205826 649454
rect 206062 649218 206146 649454
rect 206382 649218 206414 649454
rect 205794 649134 206414 649218
rect 205794 648898 205826 649134
rect 206062 648898 206146 649134
rect 206382 648898 206414 649134
rect 205794 615454 206414 648898
rect 205794 615218 205826 615454
rect 206062 615218 206146 615454
rect 206382 615218 206414 615454
rect 205794 615134 206414 615218
rect 205794 614898 205826 615134
rect 206062 614898 206146 615134
rect 206382 614898 206414 615134
rect 205794 581454 206414 614898
rect 205794 581218 205826 581454
rect 206062 581218 206146 581454
rect 206382 581218 206414 581454
rect 205794 581134 206414 581218
rect 205794 580898 205826 581134
rect 206062 580898 206146 581134
rect 206382 580898 206414 581134
rect 205794 547454 206414 580898
rect 205794 547218 205826 547454
rect 206062 547218 206146 547454
rect 206382 547218 206414 547454
rect 205794 547134 206414 547218
rect 205794 546898 205826 547134
rect 206062 546898 206146 547134
rect 206382 546898 206414 547134
rect 205794 513454 206414 546898
rect 205794 513218 205826 513454
rect 206062 513218 206146 513454
rect 206382 513218 206414 513454
rect 205794 513134 206414 513218
rect 205794 512898 205826 513134
rect 206062 512898 206146 513134
rect 206382 512898 206414 513134
rect 205794 479454 206414 512898
rect 205794 479218 205826 479454
rect 206062 479218 206146 479454
rect 206382 479218 206414 479454
rect 205794 479134 206414 479218
rect 205794 478898 205826 479134
rect 206062 478898 206146 479134
rect 206382 478898 206414 479134
rect 205794 445454 206414 478898
rect 205794 445218 205826 445454
rect 206062 445218 206146 445454
rect 206382 445218 206414 445454
rect 205794 445134 206414 445218
rect 205794 444898 205826 445134
rect 206062 444898 206146 445134
rect 206382 444898 206414 445134
rect 205794 411454 206414 444898
rect 205794 411218 205826 411454
rect 206062 411218 206146 411454
rect 206382 411218 206414 411454
rect 205794 411134 206414 411218
rect 205794 410898 205826 411134
rect 206062 410898 206146 411134
rect 206382 410898 206414 411134
rect 205794 377454 206414 410898
rect 205794 377218 205826 377454
rect 206062 377218 206146 377454
rect 206382 377218 206414 377454
rect 205794 377134 206414 377218
rect 205794 376898 205826 377134
rect 206062 376898 206146 377134
rect 206382 376898 206414 377134
rect 205794 343454 206414 376898
rect 205794 343218 205826 343454
rect 206062 343218 206146 343454
rect 206382 343218 206414 343454
rect 205794 343134 206414 343218
rect 205794 342898 205826 343134
rect 206062 342898 206146 343134
rect 206382 342898 206414 343134
rect 205794 309454 206414 342898
rect 205794 309218 205826 309454
rect 206062 309218 206146 309454
rect 206382 309218 206414 309454
rect 205794 309134 206414 309218
rect 205794 308898 205826 309134
rect 206062 308898 206146 309134
rect 206382 308898 206414 309134
rect 205794 275454 206414 308898
rect 205794 275218 205826 275454
rect 206062 275218 206146 275454
rect 206382 275218 206414 275454
rect 205794 275134 206414 275218
rect 205794 274898 205826 275134
rect 206062 274898 206146 275134
rect 206382 274898 206414 275134
rect 205794 241454 206414 274898
rect 205794 241218 205826 241454
rect 206062 241218 206146 241454
rect 206382 241218 206414 241454
rect 205794 241134 206414 241218
rect 205794 240898 205826 241134
rect 206062 240898 206146 241134
rect 206382 240898 206414 241134
rect 205794 225660 206414 240898
rect 209514 705798 210134 711590
rect 209514 705562 209546 705798
rect 209782 705562 209866 705798
rect 210102 705562 210134 705798
rect 209514 705478 210134 705562
rect 209514 705242 209546 705478
rect 209782 705242 209866 705478
rect 210102 705242 210134 705478
rect 209514 687174 210134 705242
rect 209514 686938 209546 687174
rect 209782 686938 209866 687174
rect 210102 686938 210134 687174
rect 209514 686854 210134 686938
rect 209514 686618 209546 686854
rect 209782 686618 209866 686854
rect 210102 686618 210134 686854
rect 209514 653174 210134 686618
rect 209514 652938 209546 653174
rect 209782 652938 209866 653174
rect 210102 652938 210134 653174
rect 209514 652854 210134 652938
rect 209514 652618 209546 652854
rect 209782 652618 209866 652854
rect 210102 652618 210134 652854
rect 209514 619174 210134 652618
rect 209514 618938 209546 619174
rect 209782 618938 209866 619174
rect 210102 618938 210134 619174
rect 209514 618854 210134 618938
rect 209514 618618 209546 618854
rect 209782 618618 209866 618854
rect 210102 618618 210134 618854
rect 209514 585174 210134 618618
rect 209514 584938 209546 585174
rect 209782 584938 209866 585174
rect 210102 584938 210134 585174
rect 209514 584854 210134 584938
rect 209514 584618 209546 584854
rect 209782 584618 209866 584854
rect 210102 584618 210134 584854
rect 209514 551174 210134 584618
rect 209514 550938 209546 551174
rect 209782 550938 209866 551174
rect 210102 550938 210134 551174
rect 209514 550854 210134 550938
rect 209514 550618 209546 550854
rect 209782 550618 209866 550854
rect 210102 550618 210134 550854
rect 209514 517174 210134 550618
rect 209514 516938 209546 517174
rect 209782 516938 209866 517174
rect 210102 516938 210134 517174
rect 209514 516854 210134 516938
rect 209514 516618 209546 516854
rect 209782 516618 209866 516854
rect 210102 516618 210134 516854
rect 209514 483174 210134 516618
rect 209514 482938 209546 483174
rect 209782 482938 209866 483174
rect 210102 482938 210134 483174
rect 209514 482854 210134 482938
rect 209514 482618 209546 482854
rect 209782 482618 209866 482854
rect 210102 482618 210134 482854
rect 209514 449174 210134 482618
rect 209514 448938 209546 449174
rect 209782 448938 209866 449174
rect 210102 448938 210134 449174
rect 209514 448854 210134 448938
rect 209514 448618 209546 448854
rect 209782 448618 209866 448854
rect 210102 448618 210134 448854
rect 209514 415174 210134 448618
rect 209514 414938 209546 415174
rect 209782 414938 209866 415174
rect 210102 414938 210134 415174
rect 209514 414854 210134 414938
rect 209514 414618 209546 414854
rect 209782 414618 209866 414854
rect 210102 414618 210134 414854
rect 209514 381174 210134 414618
rect 209514 380938 209546 381174
rect 209782 380938 209866 381174
rect 210102 380938 210134 381174
rect 209514 380854 210134 380938
rect 209514 380618 209546 380854
rect 209782 380618 209866 380854
rect 210102 380618 210134 380854
rect 209514 347174 210134 380618
rect 209514 346938 209546 347174
rect 209782 346938 209866 347174
rect 210102 346938 210134 347174
rect 209514 346854 210134 346938
rect 209514 346618 209546 346854
rect 209782 346618 209866 346854
rect 210102 346618 210134 346854
rect 209514 313174 210134 346618
rect 209514 312938 209546 313174
rect 209782 312938 209866 313174
rect 210102 312938 210134 313174
rect 209514 312854 210134 312938
rect 209514 312618 209546 312854
rect 209782 312618 209866 312854
rect 210102 312618 210134 312854
rect 209514 279174 210134 312618
rect 209514 278938 209546 279174
rect 209782 278938 209866 279174
rect 210102 278938 210134 279174
rect 209514 278854 210134 278938
rect 209514 278618 209546 278854
rect 209782 278618 209866 278854
rect 210102 278618 210134 278854
rect 209514 245174 210134 278618
rect 209514 244938 209546 245174
rect 209782 244938 209866 245174
rect 210102 244938 210134 245174
rect 209514 244854 210134 244938
rect 209514 244618 209546 244854
rect 209782 244618 209866 244854
rect 210102 244618 210134 244854
rect 209514 225660 210134 244618
rect 213234 706758 213854 711590
rect 213234 706522 213266 706758
rect 213502 706522 213586 706758
rect 213822 706522 213854 706758
rect 213234 706438 213854 706522
rect 213234 706202 213266 706438
rect 213502 706202 213586 706438
rect 213822 706202 213854 706438
rect 213234 690894 213854 706202
rect 213234 690658 213266 690894
rect 213502 690658 213586 690894
rect 213822 690658 213854 690894
rect 213234 690574 213854 690658
rect 213234 690338 213266 690574
rect 213502 690338 213586 690574
rect 213822 690338 213854 690574
rect 213234 656894 213854 690338
rect 213234 656658 213266 656894
rect 213502 656658 213586 656894
rect 213822 656658 213854 656894
rect 213234 656574 213854 656658
rect 213234 656338 213266 656574
rect 213502 656338 213586 656574
rect 213822 656338 213854 656574
rect 213234 622894 213854 656338
rect 213234 622658 213266 622894
rect 213502 622658 213586 622894
rect 213822 622658 213854 622894
rect 213234 622574 213854 622658
rect 213234 622338 213266 622574
rect 213502 622338 213586 622574
rect 213822 622338 213854 622574
rect 213234 588894 213854 622338
rect 213234 588658 213266 588894
rect 213502 588658 213586 588894
rect 213822 588658 213854 588894
rect 213234 588574 213854 588658
rect 213234 588338 213266 588574
rect 213502 588338 213586 588574
rect 213822 588338 213854 588574
rect 213234 554894 213854 588338
rect 213234 554658 213266 554894
rect 213502 554658 213586 554894
rect 213822 554658 213854 554894
rect 213234 554574 213854 554658
rect 213234 554338 213266 554574
rect 213502 554338 213586 554574
rect 213822 554338 213854 554574
rect 213234 520894 213854 554338
rect 213234 520658 213266 520894
rect 213502 520658 213586 520894
rect 213822 520658 213854 520894
rect 213234 520574 213854 520658
rect 213234 520338 213266 520574
rect 213502 520338 213586 520574
rect 213822 520338 213854 520574
rect 213234 486894 213854 520338
rect 213234 486658 213266 486894
rect 213502 486658 213586 486894
rect 213822 486658 213854 486894
rect 213234 486574 213854 486658
rect 213234 486338 213266 486574
rect 213502 486338 213586 486574
rect 213822 486338 213854 486574
rect 213234 452894 213854 486338
rect 213234 452658 213266 452894
rect 213502 452658 213586 452894
rect 213822 452658 213854 452894
rect 213234 452574 213854 452658
rect 213234 452338 213266 452574
rect 213502 452338 213586 452574
rect 213822 452338 213854 452574
rect 213234 418894 213854 452338
rect 213234 418658 213266 418894
rect 213502 418658 213586 418894
rect 213822 418658 213854 418894
rect 213234 418574 213854 418658
rect 213234 418338 213266 418574
rect 213502 418338 213586 418574
rect 213822 418338 213854 418574
rect 213234 384894 213854 418338
rect 213234 384658 213266 384894
rect 213502 384658 213586 384894
rect 213822 384658 213854 384894
rect 213234 384574 213854 384658
rect 213234 384338 213266 384574
rect 213502 384338 213586 384574
rect 213822 384338 213854 384574
rect 213234 350894 213854 384338
rect 213234 350658 213266 350894
rect 213502 350658 213586 350894
rect 213822 350658 213854 350894
rect 213234 350574 213854 350658
rect 213234 350338 213266 350574
rect 213502 350338 213586 350574
rect 213822 350338 213854 350574
rect 213234 316894 213854 350338
rect 213234 316658 213266 316894
rect 213502 316658 213586 316894
rect 213822 316658 213854 316894
rect 213234 316574 213854 316658
rect 213234 316338 213266 316574
rect 213502 316338 213586 316574
rect 213822 316338 213854 316574
rect 213234 282894 213854 316338
rect 213234 282658 213266 282894
rect 213502 282658 213586 282894
rect 213822 282658 213854 282894
rect 213234 282574 213854 282658
rect 213234 282338 213266 282574
rect 213502 282338 213586 282574
rect 213822 282338 213854 282574
rect 213234 248894 213854 282338
rect 213234 248658 213266 248894
rect 213502 248658 213586 248894
rect 213822 248658 213854 248894
rect 213234 248574 213854 248658
rect 213234 248338 213266 248574
rect 213502 248338 213586 248574
rect 213822 248338 213854 248574
rect 213234 225660 213854 248338
rect 216954 707718 217574 711590
rect 216954 707482 216986 707718
rect 217222 707482 217306 707718
rect 217542 707482 217574 707718
rect 216954 707398 217574 707482
rect 216954 707162 216986 707398
rect 217222 707162 217306 707398
rect 217542 707162 217574 707398
rect 216954 694614 217574 707162
rect 216954 694378 216986 694614
rect 217222 694378 217306 694614
rect 217542 694378 217574 694614
rect 216954 694294 217574 694378
rect 216954 694058 216986 694294
rect 217222 694058 217306 694294
rect 217542 694058 217574 694294
rect 216954 660614 217574 694058
rect 216954 660378 216986 660614
rect 217222 660378 217306 660614
rect 217542 660378 217574 660614
rect 216954 660294 217574 660378
rect 216954 660058 216986 660294
rect 217222 660058 217306 660294
rect 217542 660058 217574 660294
rect 216954 626614 217574 660058
rect 216954 626378 216986 626614
rect 217222 626378 217306 626614
rect 217542 626378 217574 626614
rect 216954 626294 217574 626378
rect 216954 626058 216986 626294
rect 217222 626058 217306 626294
rect 217542 626058 217574 626294
rect 216954 592614 217574 626058
rect 216954 592378 216986 592614
rect 217222 592378 217306 592614
rect 217542 592378 217574 592614
rect 216954 592294 217574 592378
rect 216954 592058 216986 592294
rect 217222 592058 217306 592294
rect 217542 592058 217574 592294
rect 216954 558614 217574 592058
rect 216954 558378 216986 558614
rect 217222 558378 217306 558614
rect 217542 558378 217574 558614
rect 216954 558294 217574 558378
rect 216954 558058 216986 558294
rect 217222 558058 217306 558294
rect 217542 558058 217574 558294
rect 216954 524614 217574 558058
rect 216954 524378 216986 524614
rect 217222 524378 217306 524614
rect 217542 524378 217574 524614
rect 216954 524294 217574 524378
rect 216954 524058 216986 524294
rect 217222 524058 217306 524294
rect 217542 524058 217574 524294
rect 216954 490614 217574 524058
rect 216954 490378 216986 490614
rect 217222 490378 217306 490614
rect 217542 490378 217574 490614
rect 216954 490294 217574 490378
rect 216954 490058 216986 490294
rect 217222 490058 217306 490294
rect 217542 490058 217574 490294
rect 216954 456614 217574 490058
rect 216954 456378 216986 456614
rect 217222 456378 217306 456614
rect 217542 456378 217574 456614
rect 216954 456294 217574 456378
rect 216954 456058 216986 456294
rect 217222 456058 217306 456294
rect 217542 456058 217574 456294
rect 216954 422614 217574 456058
rect 216954 422378 216986 422614
rect 217222 422378 217306 422614
rect 217542 422378 217574 422614
rect 216954 422294 217574 422378
rect 216954 422058 216986 422294
rect 217222 422058 217306 422294
rect 217542 422058 217574 422294
rect 216954 388614 217574 422058
rect 216954 388378 216986 388614
rect 217222 388378 217306 388614
rect 217542 388378 217574 388614
rect 216954 388294 217574 388378
rect 216954 388058 216986 388294
rect 217222 388058 217306 388294
rect 217542 388058 217574 388294
rect 216954 354614 217574 388058
rect 216954 354378 216986 354614
rect 217222 354378 217306 354614
rect 217542 354378 217574 354614
rect 216954 354294 217574 354378
rect 216954 354058 216986 354294
rect 217222 354058 217306 354294
rect 217542 354058 217574 354294
rect 216954 320614 217574 354058
rect 216954 320378 216986 320614
rect 217222 320378 217306 320614
rect 217542 320378 217574 320614
rect 216954 320294 217574 320378
rect 216954 320058 216986 320294
rect 217222 320058 217306 320294
rect 217542 320058 217574 320294
rect 216954 286614 217574 320058
rect 216954 286378 216986 286614
rect 217222 286378 217306 286614
rect 217542 286378 217574 286614
rect 216954 286294 217574 286378
rect 216954 286058 216986 286294
rect 217222 286058 217306 286294
rect 217542 286058 217574 286294
rect 216954 252614 217574 286058
rect 216954 252378 216986 252614
rect 217222 252378 217306 252614
rect 217542 252378 217574 252614
rect 216954 252294 217574 252378
rect 216954 252058 216986 252294
rect 217222 252058 217306 252294
rect 217542 252058 217574 252294
rect 216954 225660 217574 252058
rect 220674 708678 221294 711590
rect 220674 708442 220706 708678
rect 220942 708442 221026 708678
rect 221262 708442 221294 708678
rect 220674 708358 221294 708442
rect 220674 708122 220706 708358
rect 220942 708122 221026 708358
rect 221262 708122 221294 708358
rect 220674 698334 221294 708122
rect 220674 698098 220706 698334
rect 220942 698098 221026 698334
rect 221262 698098 221294 698334
rect 220674 698014 221294 698098
rect 220674 697778 220706 698014
rect 220942 697778 221026 698014
rect 221262 697778 221294 698014
rect 220674 664334 221294 697778
rect 220674 664098 220706 664334
rect 220942 664098 221026 664334
rect 221262 664098 221294 664334
rect 220674 664014 221294 664098
rect 220674 663778 220706 664014
rect 220942 663778 221026 664014
rect 221262 663778 221294 664014
rect 220674 630334 221294 663778
rect 220674 630098 220706 630334
rect 220942 630098 221026 630334
rect 221262 630098 221294 630334
rect 220674 630014 221294 630098
rect 220674 629778 220706 630014
rect 220942 629778 221026 630014
rect 221262 629778 221294 630014
rect 220674 596334 221294 629778
rect 220674 596098 220706 596334
rect 220942 596098 221026 596334
rect 221262 596098 221294 596334
rect 220674 596014 221294 596098
rect 220674 595778 220706 596014
rect 220942 595778 221026 596014
rect 221262 595778 221294 596014
rect 220674 562334 221294 595778
rect 220674 562098 220706 562334
rect 220942 562098 221026 562334
rect 221262 562098 221294 562334
rect 220674 562014 221294 562098
rect 220674 561778 220706 562014
rect 220942 561778 221026 562014
rect 221262 561778 221294 562014
rect 220674 528334 221294 561778
rect 220674 528098 220706 528334
rect 220942 528098 221026 528334
rect 221262 528098 221294 528334
rect 220674 528014 221294 528098
rect 220674 527778 220706 528014
rect 220942 527778 221026 528014
rect 221262 527778 221294 528014
rect 220674 494334 221294 527778
rect 220674 494098 220706 494334
rect 220942 494098 221026 494334
rect 221262 494098 221294 494334
rect 220674 494014 221294 494098
rect 220674 493778 220706 494014
rect 220942 493778 221026 494014
rect 221262 493778 221294 494014
rect 220674 460334 221294 493778
rect 220674 460098 220706 460334
rect 220942 460098 221026 460334
rect 221262 460098 221294 460334
rect 220674 460014 221294 460098
rect 220674 459778 220706 460014
rect 220942 459778 221026 460014
rect 221262 459778 221294 460014
rect 220674 426334 221294 459778
rect 220674 426098 220706 426334
rect 220942 426098 221026 426334
rect 221262 426098 221294 426334
rect 220674 426014 221294 426098
rect 220674 425778 220706 426014
rect 220942 425778 221026 426014
rect 221262 425778 221294 426014
rect 220674 392334 221294 425778
rect 220674 392098 220706 392334
rect 220942 392098 221026 392334
rect 221262 392098 221294 392334
rect 220674 392014 221294 392098
rect 220674 391778 220706 392014
rect 220942 391778 221026 392014
rect 221262 391778 221294 392014
rect 220674 358334 221294 391778
rect 220674 358098 220706 358334
rect 220942 358098 221026 358334
rect 221262 358098 221294 358334
rect 220674 358014 221294 358098
rect 220674 357778 220706 358014
rect 220942 357778 221026 358014
rect 221262 357778 221294 358014
rect 220674 324334 221294 357778
rect 220674 324098 220706 324334
rect 220942 324098 221026 324334
rect 221262 324098 221294 324334
rect 220674 324014 221294 324098
rect 220674 323778 220706 324014
rect 220942 323778 221026 324014
rect 221262 323778 221294 324014
rect 220674 290334 221294 323778
rect 220674 290098 220706 290334
rect 220942 290098 221026 290334
rect 221262 290098 221294 290334
rect 220674 290014 221294 290098
rect 220674 289778 220706 290014
rect 220942 289778 221026 290014
rect 221262 289778 221294 290014
rect 220674 256334 221294 289778
rect 220674 256098 220706 256334
rect 220942 256098 221026 256334
rect 221262 256098 221294 256334
rect 220674 256014 221294 256098
rect 220674 255778 220706 256014
rect 220942 255778 221026 256014
rect 221262 255778 221294 256014
rect 160114 195538 160146 195774
rect 160382 195538 160466 195774
rect 160702 195538 160734 195774
rect 160114 195454 160734 195538
rect 160114 195218 160146 195454
rect 160382 195218 160466 195454
rect 160702 195218 160734 195454
rect 160114 194880 160734 195218
rect 163834 199494 164454 214340
rect 163834 199258 163866 199494
rect 164102 199258 164186 199494
rect 164422 199258 164454 199494
rect 163834 199174 164454 199258
rect 163834 198938 163866 199174
rect 164102 198938 164186 199174
rect 164422 198938 164454 199174
rect 134314 188334 162514 188366
rect 134314 188098 134376 188334
rect 134612 188098 134696 188334
rect 134932 188098 135016 188334
rect 135252 188098 135336 188334
rect 135572 188098 135656 188334
rect 135892 188098 135976 188334
rect 136212 188098 136296 188334
rect 136532 188098 136616 188334
rect 136852 188098 136936 188334
rect 137172 188098 137256 188334
rect 137492 188098 137576 188334
rect 137812 188098 137896 188334
rect 138132 188098 138216 188334
rect 138452 188098 138536 188334
rect 138772 188098 138856 188334
rect 139092 188098 139176 188334
rect 139412 188098 139496 188334
rect 139732 188098 139816 188334
rect 140052 188098 140136 188334
rect 140372 188098 140456 188334
rect 140692 188098 140776 188334
rect 141012 188098 141096 188334
rect 141332 188098 141416 188334
rect 141652 188098 141736 188334
rect 141972 188098 142056 188334
rect 142292 188098 142376 188334
rect 142612 188098 142696 188334
rect 142932 188098 143016 188334
rect 143252 188098 143336 188334
rect 143572 188098 143656 188334
rect 143892 188098 143976 188334
rect 144212 188098 144296 188334
rect 144532 188098 144616 188334
rect 144852 188098 144936 188334
rect 145172 188098 145256 188334
rect 145492 188098 145576 188334
rect 145812 188098 145896 188334
rect 146132 188098 146216 188334
rect 146452 188098 146536 188334
rect 146772 188098 146856 188334
rect 147092 188098 147176 188334
rect 147412 188098 147496 188334
rect 147732 188098 147816 188334
rect 148052 188098 148136 188334
rect 148372 188098 148456 188334
rect 148692 188098 148776 188334
rect 149012 188098 149096 188334
rect 149332 188098 149416 188334
rect 149652 188098 149736 188334
rect 149972 188098 150056 188334
rect 150292 188098 150376 188334
rect 150612 188098 150696 188334
rect 150932 188098 151016 188334
rect 151252 188098 151336 188334
rect 151572 188098 151656 188334
rect 151892 188098 151976 188334
rect 152212 188098 152296 188334
rect 152532 188098 152616 188334
rect 152852 188098 152936 188334
rect 153172 188098 153256 188334
rect 153492 188098 153576 188334
rect 153812 188098 153896 188334
rect 154132 188098 154216 188334
rect 154452 188098 154536 188334
rect 154772 188098 154856 188334
rect 155092 188098 155176 188334
rect 155412 188098 155496 188334
rect 155732 188098 155816 188334
rect 156052 188098 156136 188334
rect 156372 188098 156456 188334
rect 156692 188098 156776 188334
rect 157012 188098 157096 188334
rect 157332 188098 157416 188334
rect 157652 188098 157736 188334
rect 157972 188098 158056 188334
rect 158292 188098 158376 188334
rect 158612 188098 158696 188334
rect 158932 188098 159016 188334
rect 159252 188098 159336 188334
rect 159572 188098 159656 188334
rect 159892 188098 159976 188334
rect 160212 188098 160296 188334
rect 160532 188098 160616 188334
rect 160852 188098 160936 188334
rect 161172 188098 161256 188334
rect 161492 188098 161576 188334
rect 161812 188098 161896 188334
rect 162132 188098 162216 188334
rect 162452 188098 162514 188334
rect 134314 188014 162514 188098
rect 134314 187778 134376 188014
rect 134612 187778 134696 188014
rect 134932 187778 135016 188014
rect 135252 187778 135336 188014
rect 135572 187778 135656 188014
rect 135892 187778 135976 188014
rect 136212 187778 136296 188014
rect 136532 187778 136616 188014
rect 136852 187778 136936 188014
rect 137172 187778 137256 188014
rect 137492 187778 137576 188014
rect 137812 187778 137896 188014
rect 138132 187778 138216 188014
rect 138452 187778 138536 188014
rect 138772 187778 138856 188014
rect 139092 187778 139176 188014
rect 139412 187778 139496 188014
rect 139732 187778 139816 188014
rect 140052 187778 140136 188014
rect 140372 187778 140456 188014
rect 140692 187778 140776 188014
rect 141012 187778 141096 188014
rect 141332 187778 141416 188014
rect 141652 187778 141736 188014
rect 141972 187778 142056 188014
rect 142292 187778 142376 188014
rect 142612 187778 142696 188014
rect 142932 187778 143016 188014
rect 143252 187778 143336 188014
rect 143572 187778 143656 188014
rect 143892 187778 143976 188014
rect 144212 187778 144296 188014
rect 144532 187778 144616 188014
rect 144852 187778 144936 188014
rect 145172 187778 145256 188014
rect 145492 187778 145576 188014
rect 145812 187778 145896 188014
rect 146132 187778 146216 188014
rect 146452 187778 146536 188014
rect 146772 187778 146856 188014
rect 147092 187778 147176 188014
rect 147412 187778 147496 188014
rect 147732 187778 147816 188014
rect 148052 187778 148136 188014
rect 148372 187778 148456 188014
rect 148692 187778 148776 188014
rect 149012 187778 149096 188014
rect 149332 187778 149416 188014
rect 149652 187778 149736 188014
rect 149972 187778 150056 188014
rect 150292 187778 150376 188014
rect 150612 187778 150696 188014
rect 150932 187778 151016 188014
rect 151252 187778 151336 188014
rect 151572 187778 151656 188014
rect 151892 187778 151976 188014
rect 152212 187778 152296 188014
rect 152532 187778 152616 188014
rect 152852 187778 152936 188014
rect 153172 187778 153256 188014
rect 153492 187778 153576 188014
rect 153812 187778 153896 188014
rect 154132 187778 154216 188014
rect 154452 187778 154536 188014
rect 154772 187778 154856 188014
rect 155092 187778 155176 188014
rect 155412 187778 155496 188014
rect 155732 187778 155816 188014
rect 156052 187778 156136 188014
rect 156372 187778 156456 188014
rect 156692 187778 156776 188014
rect 157012 187778 157096 188014
rect 157332 187778 157416 188014
rect 157652 187778 157736 188014
rect 157972 187778 158056 188014
rect 158292 187778 158376 188014
rect 158612 187778 158696 188014
rect 158932 187778 159016 188014
rect 159252 187778 159336 188014
rect 159572 187778 159656 188014
rect 159892 187778 159976 188014
rect 160212 187778 160296 188014
rect 160532 187778 160616 188014
rect 160852 187778 160936 188014
rect 161172 187778 161256 188014
rect 161492 187778 161576 188014
rect 161812 187778 161896 188014
rect 162132 187778 162216 188014
rect 162452 187778 162514 188014
rect 134314 187746 162514 187778
rect 136035 181116 136101 181117
rect 136035 181052 136036 181116
rect 136100 181052 136101 181116
rect 136035 181051 136101 181052
rect 135851 180980 135917 180981
rect 135851 180916 135852 180980
rect 135916 180916 135917 180980
rect 135851 180915 135917 180916
rect 129834 165258 129866 165494
rect 130102 165258 130186 165494
rect 130422 165258 130454 165494
rect 129834 165174 130454 165258
rect 129834 164938 129866 165174
rect 130102 164938 130186 165174
rect 130422 164938 130454 165174
rect 129834 134417 130454 164938
rect 134414 161781 135034 161806
rect 134414 161545 134446 161781
rect 134682 161545 134766 161781
rect 135002 161545 135034 161781
rect 134414 161461 135034 161545
rect 135854 161533 135914 180915
rect 136038 171150 136098 181051
rect 137794 173454 138414 185520
rect 145234 180894 145854 185520
rect 145234 180658 145266 180894
rect 145502 180658 145586 180894
rect 145822 180658 145854 180894
rect 145234 180574 145854 180658
rect 145234 180338 145266 180574
rect 145502 180338 145586 180574
rect 145822 180338 145854 180574
rect 145234 179075 145854 180338
rect 148954 184614 149574 185520
rect 148954 184378 148986 184614
rect 149222 184378 149306 184614
rect 149542 184378 149574 184614
rect 148954 184294 149574 184378
rect 148954 184058 148986 184294
rect 149222 184058 149306 184294
rect 149542 184058 149574 184294
rect 148954 179075 149574 184058
rect 140635 178132 140701 178133
rect 140635 178068 140636 178132
rect 140700 178068 140701 178132
rect 140635 178067 140701 178068
rect 139531 177444 139597 177445
rect 139531 177380 139532 177444
rect 139596 177380 139597 177444
rect 139531 177379 139597 177380
rect 137794 173218 137826 173454
rect 138062 173218 138146 173454
rect 138382 173218 138414 173454
rect 137794 173134 138414 173218
rect 137794 172898 137826 173134
rect 138062 172898 138146 173134
rect 138382 172898 138414 173134
rect 136038 171090 136466 171150
rect 135851 161532 135917 161533
rect 135851 161468 135852 161532
rect 135916 161468 135917 161532
rect 135851 161467 135917 161468
rect 134414 161225 134446 161461
rect 134682 161225 134766 161461
rect 135002 161225 135034 161461
rect 136406 161397 136466 171090
rect 137794 163280 138414 172898
rect 139534 165205 139594 177379
rect 139531 165204 139597 165205
rect 139531 165140 139532 165204
rect 139596 165140 139597 165204
rect 139531 165139 139597 165140
rect 136403 161396 136469 161397
rect 136403 161332 136404 161396
rect 136468 161332 136469 161396
rect 136403 161331 136469 161332
rect 134414 161200 135034 161225
rect 135851 160036 135917 160037
rect 135851 159972 135852 160036
rect 135916 159972 135917 160036
rect 135851 159971 135917 159972
rect 136035 160036 136101 160037
rect 136035 159972 136036 160036
rect 136100 159972 136101 160036
rect 136035 159971 136101 159972
rect 135854 137597 135914 159971
rect 135851 137596 135917 137597
rect 135851 137532 135852 137596
rect 135916 137532 135917 137596
rect 135851 137531 135917 137532
rect 136038 137461 136098 159971
rect 140638 152421 140698 178067
rect 141923 176084 141989 176085
rect 141923 176020 141924 176084
rect 141988 176020 141989 176084
rect 141923 176019 141989 176020
rect 141555 172548 141621 172549
rect 141555 172484 141556 172548
rect 141620 172484 141621 172548
rect 141555 172483 141621 172484
rect 141558 162213 141618 172483
rect 141555 162212 141621 162213
rect 141555 162148 141556 162212
rect 141620 162148 141621 162212
rect 141555 162147 141621 162148
rect 140635 152420 140701 152421
rect 140635 152356 140636 152420
rect 140700 152356 140701 152420
rect 140635 152355 140701 152356
rect 141926 137461 141986 176019
rect 160114 161774 160734 165832
rect 160114 161538 160146 161774
rect 160382 161538 160466 161774
rect 160702 161538 160734 161774
rect 160114 161454 160734 161538
rect 160114 161218 160146 161454
rect 160382 161218 160466 161454
rect 160702 161218 160734 161454
rect 136035 137460 136101 137461
rect 136035 137396 136036 137460
rect 136100 137396 136101 137460
rect 136035 137395 136101 137396
rect 141923 137460 141989 137461
rect 141923 137396 141924 137460
rect 141988 137396 141989 137460
rect 141923 137395 141989 137396
rect 160114 134417 160734 161218
rect 163834 165494 164454 198938
rect 163834 165258 163866 165494
rect 164102 165258 164186 165494
rect 164422 165258 164454 165494
rect 163834 165174 164454 165258
rect 163834 164938 163866 165174
rect 164102 164938 164186 165174
rect 164422 164938 164454 165174
rect 163834 134417 164454 164938
rect 171794 207454 172414 214340
rect 171794 207218 171826 207454
rect 172062 207218 172146 207454
rect 172382 207218 172414 207454
rect 171794 207134 172414 207218
rect 171794 206898 171826 207134
rect 172062 206898 172146 207134
rect 172382 206898 172414 207134
rect 171794 173454 172414 206898
rect 171794 173218 171826 173454
rect 172062 173218 172146 173454
rect 172382 173218 172414 173454
rect 171794 173134 172414 173218
rect 171794 172898 171826 173134
rect 172062 172898 172146 173134
rect 172382 172898 172414 173134
rect 171794 139454 172414 172898
rect 171794 139218 171826 139454
rect 172062 139218 172146 139454
rect 172382 139218 172414 139454
rect 171794 139134 172414 139218
rect 171794 138898 171826 139134
rect 172062 138898 172146 139134
rect 172382 138898 172414 139134
rect 114954 116378 114986 116614
rect 115222 116378 115306 116614
rect 115542 116378 115574 116614
rect 114954 116294 115574 116378
rect 114954 116058 114986 116294
rect 115222 116058 115306 116294
rect 115542 116058 115574 116294
rect 114954 82614 115574 116058
rect 135568 109174 135888 109206
rect 135568 108938 135610 109174
rect 135846 108938 135888 109174
rect 135568 108854 135888 108938
rect 135568 108618 135610 108854
rect 135846 108618 135888 108854
rect 135568 108586 135888 108618
rect 166288 109174 166608 109206
rect 166288 108938 166330 109174
rect 166566 108938 166608 109174
rect 166288 108854 166608 108938
rect 166288 108618 166330 108854
rect 166566 108618 166608 108854
rect 166288 108586 166608 108618
rect 120208 105454 120528 105486
rect 120208 105218 120250 105454
rect 120486 105218 120528 105454
rect 120208 105134 120528 105218
rect 120208 104898 120250 105134
rect 120486 104898 120528 105134
rect 120208 104866 120528 104898
rect 150928 105454 151248 105486
rect 150928 105218 150970 105454
rect 151206 105218 151248 105454
rect 150928 105134 151248 105218
rect 150928 104898 150970 105134
rect 151206 104898 151248 105134
rect 150928 104866 151248 104898
rect 171794 105454 172414 138898
rect 171794 105218 171826 105454
rect 172062 105218 172146 105454
rect 172382 105218 172414 105454
rect 171794 105134 172414 105218
rect 171794 104898 171826 105134
rect 172062 104898 172146 105134
rect 172382 104898 172414 105134
rect 114954 82378 114986 82614
rect 115222 82378 115306 82614
rect 115542 82378 115574 82614
rect 114954 82294 115574 82378
rect 114954 82058 114986 82294
rect 115222 82058 115306 82294
rect 115542 82058 115574 82294
rect 114954 48614 115574 82058
rect 169339 75444 169405 75445
rect 169339 75380 169340 75444
rect 169404 75380 169405 75444
rect 169339 75379 169405 75380
rect 147443 75308 147509 75309
rect 147443 75244 147444 75308
rect 147508 75244 147509 75308
rect 147443 75243 147509 75244
rect 114954 48378 114986 48614
rect 115222 48378 115306 48614
rect 115542 48378 115574 48614
rect 114954 48294 115574 48378
rect 114954 48058 114986 48294
rect 115222 48058 115306 48294
rect 115542 48058 115574 48294
rect 114954 14614 115574 48058
rect 114954 14378 114986 14614
rect 115222 14378 115306 14614
rect 115542 14378 115574 14614
rect 114954 14294 115574 14378
rect 114954 14058 114986 14294
rect 115222 14058 115306 14294
rect 115542 14058 115574 14294
rect 114954 -3226 115574 14058
rect 114954 -3462 114986 -3226
rect 115222 -3462 115306 -3226
rect 115542 -3462 115574 -3226
rect 114954 -3546 115574 -3462
rect 114954 -3782 114986 -3546
rect 115222 -3782 115306 -3546
rect 115542 -3782 115574 -3546
rect 114954 -7654 115574 -3782
rect 118674 52334 119294 74063
rect 121499 72724 121565 72725
rect 121499 72660 121500 72724
rect 121564 72660 121565 72724
rect 121499 72659 121565 72660
rect 121502 69597 121562 72659
rect 121499 69596 121565 69597
rect 121499 69532 121500 69596
rect 121564 69532 121565 69596
rect 121499 69531 121565 69532
rect 118674 52098 118706 52334
rect 118942 52098 119026 52334
rect 119262 52098 119294 52334
rect 118674 52014 119294 52098
rect 118674 51778 118706 52014
rect 118942 51778 119026 52014
rect 119262 51778 119294 52014
rect 118674 18334 119294 51778
rect 118674 18098 118706 18334
rect 118942 18098 119026 18334
rect 119262 18098 119294 18334
rect 118674 18014 119294 18098
rect 118674 17778 118706 18014
rect 118942 17778 119026 18014
rect 119262 17778 119294 18014
rect 118674 -4186 119294 17778
rect 118674 -4422 118706 -4186
rect 118942 -4422 119026 -4186
rect 119262 -4422 119294 -4186
rect 118674 -4506 119294 -4422
rect 118674 -4742 118706 -4506
rect 118942 -4742 119026 -4506
rect 119262 -4742 119294 -4506
rect 118674 -7654 119294 -4742
rect 122394 56054 123014 74063
rect 123707 73540 123773 73541
rect 123707 73476 123708 73540
rect 123772 73476 123773 73540
rect 123707 73475 123773 73476
rect 123155 72724 123221 72725
rect 123155 72660 123156 72724
rect 123220 72660 123221 72724
rect 123155 72659 123221 72660
rect 123158 66877 123218 72659
rect 123710 72589 123770 73475
rect 124443 72860 124509 72861
rect 124443 72796 124444 72860
rect 124508 72796 124509 72860
rect 124443 72795 124509 72796
rect 125547 72860 125613 72861
rect 125547 72796 125548 72860
rect 125612 72796 125613 72860
rect 125547 72795 125613 72796
rect 124259 72724 124325 72725
rect 124259 72660 124260 72724
rect 124324 72660 124325 72724
rect 124259 72659 124325 72660
rect 123707 72588 123773 72589
rect 123707 72524 123708 72588
rect 123772 72524 123773 72588
rect 123707 72523 123773 72524
rect 123339 72452 123405 72453
rect 123339 72388 123340 72452
rect 123404 72388 123405 72452
rect 123339 72387 123405 72388
rect 123155 66876 123221 66877
rect 123155 66812 123156 66876
rect 123220 66812 123221 66876
rect 123155 66811 123221 66812
rect 122394 55818 122426 56054
rect 122662 55818 122746 56054
rect 122982 55818 123014 56054
rect 122394 55734 123014 55818
rect 122394 55498 122426 55734
rect 122662 55498 122746 55734
rect 122982 55498 123014 55734
rect 122394 22054 123014 55498
rect 123342 51781 123402 72387
rect 124262 67013 124322 72659
rect 124259 67012 124325 67013
rect 124259 66948 124260 67012
rect 124324 66948 124325 67012
rect 124259 66947 124325 66948
rect 123339 51780 123405 51781
rect 123339 51716 123340 51780
rect 123404 51716 123405 51780
rect 123339 51715 123405 51716
rect 124446 50285 124506 72795
rect 124627 72724 124693 72725
rect 124627 72660 124628 72724
rect 124692 72660 124693 72724
rect 124627 72659 124693 72660
rect 124630 53141 124690 72659
rect 124811 72588 124877 72589
rect 124811 72524 124812 72588
rect 124876 72524 124877 72588
rect 124811 72523 124877 72524
rect 124627 53140 124693 53141
rect 124627 53076 124628 53140
rect 124692 53076 124693 53140
rect 124627 53075 124693 53076
rect 124443 50284 124509 50285
rect 124443 50220 124444 50284
rect 124508 50220 124509 50284
rect 124443 50219 124509 50220
rect 124814 48925 124874 72523
rect 124811 48924 124877 48925
rect 124811 48860 124812 48924
rect 124876 48860 124877 48924
rect 124811 48859 124877 48860
rect 125550 46205 125610 72795
rect 125731 72724 125797 72725
rect 125731 72660 125732 72724
rect 125796 72660 125797 72724
rect 125731 72659 125797 72660
rect 125734 64157 125794 72659
rect 125731 64156 125797 64157
rect 125731 64092 125732 64156
rect 125796 64092 125797 64156
rect 125731 64091 125797 64092
rect 126114 59774 126734 74063
rect 127387 72860 127453 72861
rect 127387 72796 127388 72860
rect 127452 72796 127453 72860
rect 127387 72795 127453 72796
rect 128675 72860 128741 72861
rect 128675 72796 128676 72860
rect 128740 72796 128741 72860
rect 128675 72795 128741 72796
rect 127203 72724 127269 72725
rect 127203 72660 127204 72724
rect 127268 72660 127269 72724
rect 127203 72659 127269 72660
rect 127019 72452 127085 72453
rect 127019 72388 127020 72452
rect 127084 72388 127085 72452
rect 127019 72387 127085 72388
rect 126114 59538 126146 59774
rect 126382 59538 126466 59774
rect 126702 59538 126734 59774
rect 126114 59454 126734 59538
rect 126114 59218 126146 59454
rect 126382 59218 126466 59454
rect 126702 59218 126734 59454
rect 125547 46204 125613 46205
rect 125547 46140 125548 46204
rect 125612 46140 125613 46204
rect 125547 46139 125613 46140
rect 122394 21818 122426 22054
rect 122662 21818 122746 22054
rect 122982 21818 123014 22054
rect 122394 21734 123014 21818
rect 122394 21498 122426 21734
rect 122662 21498 122746 21734
rect 122982 21498 123014 21734
rect 122394 -5146 123014 21498
rect 122394 -5382 122426 -5146
rect 122662 -5382 122746 -5146
rect 122982 -5382 123014 -5146
rect 122394 -5466 123014 -5382
rect 122394 -5702 122426 -5466
rect 122662 -5702 122746 -5466
rect 122982 -5702 123014 -5466
rect 122394 -7654 123014 -5702
rect 126114 25774 126734 59218
rect 127022 49061 127082 72387
rect 127206 50421 127266 72659
rect 127390 58717 127450 72795
rect 128491 72724 128557 72725
rect 128491 72660 128492 72724
rect 128556 72660 128557 72724
rect 128491 72659 128557 72660
rect 127571 72588 127637 72589
rect 127571 72524 127572 72588
rect 127636 72524 127637 72588
rect 127571 72523 127637 72524
rect 127574 68237 127634 72523
rect 127571 68236 127637 68237
rect 127571 68172 127572 68236
rect 127636 68172 127637 68236
rect 127571 68171 127637 68172
rect 127387 58716 127453 58717
rect 127387 58652 127388 58716
rect 127452 58652 127453 58716
rect 127387 58651 127453 58652
rect 128494 55861 128554 72659
rect 128678 61437 128738 72795
rect 128859 72588 128925 72589
rect 128859 72524 128860 72588
rect 128924 72524 128925 72588
rect 128859 72523 128925 72524
rect 128675 61436 128741 61437
rect 128675 61372 128676 61436
rect 128740 61372 128741 61436
rect 128675 61371 128741 61372
rect 128491 55860 128557 55861
rect 128491 55796 128492 55860
rect 128556 55796 128557 55860
rect 128491 55795 128557 55796
rect 127203 50420 127269 50421
rect 127203 50356 127204 50420
rect 127268 50356 127269 50420
rect 127203 50355 127269 50356
rect 127019 49060 127085 49061
rect 127019 48996 127020 49060
rect 127084 48996 127085 49060
rect 127019 48995 127085 48996
rect 126114 25538 126146 25774
rect 126382 25538 126466 25774
rect 126702 25538 126734 25774
rect 126114 25454 126734 25538
rect 126114 25218 126146 25454
rect 126382 25218 126466 25454
rect 126702 25218 126734 25454
rect 126114 -6106 126734 25218
rect 128862 6221 128922 72523
rect 129834 63494 130454 74063
rect 130883 72996 130949 72997
rect 130883 72932 130884 72996
rect 130948 72932 130949 72996
rect 130883 72931 130949 72932
rect 129834 63258 129866 63494
rect 130102 63258 130186 63494
rect 130422 63258 130454 63494
rect 129834 63174 130454 63258
rect 129834 62938 129866 63174
rect 130102 62938 130186 63174
rect 130422 62938 130454 63174
rect 129834 29494 130454 62938
rect 129834 29258 129866 29494
rect 130102 29258 130186 29494
rect 130422 29258 130454 29494
rect 129834 29174 130454 29258
rect 129834 28938 129866 29174
rect 130102 28938 130186 29174
rect 130422 28938 130454 29174
rect 128859 6220 128925 6221
rect 128859 6156 128860 6220
rect 128924 6156 128925 6220
rect 128859 6155 128925 6156
rect 126114 -6342 126146 -6106
rect 126382 -6342 126466 -6106
rect 126702 -6342 126734 -6106
rect 126114 -6426 126734 -6342
rect 126114 -6662 126146 -6426
rect 126382 -6662 126466 -6426
rect 126702 -6662 126734 -6426
rect 126114 -7654 126734 -6662
rect 129834 -7066 130454 28938
rect 130886 3909 130946 72931
rect 131987 72860 132053 72861
rect 131987 72796 131988 72860
rect 132052 72796 132053 72860
rect 131987 72795 132053 72796
rect 133275 72860 133341 72861
rect 133275 72796 133276 72860
rect 133340 72796 133341 72860
rect 133275 72795 133341 72796
rect 135115 72860 135181 72861
rect 135115 72796 135116 72860
rect 135180 72796 135181 72860
rect 135115 72795 135181 72796
rect 136587 72860 136653 72861
rect 136587 72796 136588 72860
rect 136652 72796 136653 72860
rect 136587 72795 136653 72796
rect 137323 72860 137389 72861
rect 137323 72796 137324 72860
rect 137388 72796 137389 72860
rect 137323 72795 137389 72796
rect 131990 17237 132050 72795
rect 132355 72724 132421 72725
rect 132355 72660 132356 72724
rect 132420 72660 132421 72724
rect 132355 72659 132421 72660
rect 132171 72316 132237 72317
rect 132171 72252 132172 72316
rect 132236 72252 132237 72316
rect 132171 72251 132237 72252
rect 131987 17236 132053 17237
rect 131987 17172 131988 17236
rect 132052 17172 132053 17236
rect 131987 17171 132053 17172
rect 132174 6493 132234 72251
rect 132171 6492 132237 6493
rect 132171 6428 132172 6492
rect 132236 6428 132237 6492
rect 132171 6427 132237 6428
rect 130883 3908 130949 3909
rect 130883 3844 130884 3908
rect 130948 3844 130949 3908
rect 130883 3843 130949 3844
rect 132358 3365 132418 72659
rect 133091 72588 133157 72589
rect 133091 72524 133092 72588
rect 133156 72524 133157 72588
rect 133091 72523 133157 72524
rect 133094 48245 133154 72523
rect 133091 48244 133157 48245
rect 133091 48180 133092 48244
rect 133156 48180 133157 48244
rect 133091 48179 133157 48180
rect 133278 42125 133338 72795
rect 133643 72724 133709 72725
rect 133643 72660 133644 72724
rect 133708 72660 133709 72724
rect 133643 72659 133709 72660
rect 134931 72724 134997 72725
rect 134931 72660 134932 72724
rect 134996 72660 134997 72724
rect 134931 72659 134997 72660
rect 133459 72452 133525 72453
rect 133459 72388 133460 72452
rect 133524 72388 133525 72452
rect 133459 72387 133525 72388
rect 133275 42124 133341 42125
rect 133275 42060 133276 42124
rect 133340 42060 133341 42124
rect 133275 42059 133341 42060
rect 133462 38045 133522 72387
rect 133459 38044 133525 38045
rect 133459 37980 133460 38044
rect 133524 37980 133525 38044
rect 133459 37979 133525 37980
rect 133646 15877 133706 72659
rect 134747 72588 134813 72589
rect 134747 72524 134748 72588
rect 134812 72524 134813 72588
rect 134747 72523 134813 72524
rect 134563 72452 134629 72453
rect 134563 72388 134564 72452
rect 134628 72388 134629 72452
rect 134563 72387 134629 72388
rect 134566 68645 134626 72387
rect 134563 68644 134629 68645
rect 134563 68580 134564 68644
rect 134628 68580 134629 68644
rect 134563 68579 134629 68580
rect 134750 64157 134810 72523
rect 134747 64156 134813 64157
rect 134747 64092 134748 64156
rect 134812 64092 134813 64156
rect 134747 64091 134813 64092
rect 134934 62797 134994 72659
rect 134931 62796 134997 62797
rect 134931 62732 134932 62796
rect 134996 62732 134997 62796
rect 134931 62731 134997 62732
rect 135118 52053 135178 72795
rect 136403 72724 136469 72725
rect 136403 72660 136404 72724
rect 136468 72660 136469 72724
rect 136403 72659 136469 72660
rect 136219 72588 136285 72589
rect 136219 72524 136220 72588
rect 136284 72524 136285 72588
rect 136219 72523 136285 72524
rect 136035 72452 136101 72453
rect 136035 72388 136036 72452
rect 136100 72388 136101 72452
rect 136035 72387 136101 72388
rect 136038 61437 136098 72387
rect 136035 61436 136101 61437
rect 136035 61372 136036 61436
rect 136100 61372 136101 61436
rect 136035 61371 136101 61372
rect 136222 57493 136282 72523
rect 136219 57492 136285 57493
rect 136219 57428 136220 57492
rect 136284 57428 136285 57492
rect 136219 57427 136285 57428
rect 135115 52052 135181 52053
rect 135115 51988 135116 52052
rect 135180 51988 135181 52052
rect 135115 51987 135181 51988
rect 136406 39405 136466 72659
rect 136590 68509 136650 72795
rect 136587 68508 136653 68509
rect 136587 68444 136588 68508
rect 136652 68444 136653 68508
rect 136587 68443 136653 68444
rect 137326 55997 137386 72795
rect 137507 72724 137573 72725
rect 137507 72660 137508 72724
rect 137572 72660 137573 72724
rect 137507 72659 137573 72660
rect 137323 55996 137389 55997
rect 137323 55932 137324 55996
rect 137388 55932 137389 55996
rect 137323 55931 137389 55932
rect 136403 39404 136469 39405
rect 136403 39340 136404 39404
rect 136468 39340 136469 39404
rect 136403 39339 136469 39340
rect 137510 27029 137570 72659
rect 137794 71454 138414 74063
rect 140267 73676 140333 73677
rect 140267 73612 140268 73676
rect 140332 73612 140333 73676
rect 140267 73611 140333 73612
rect 139163 73540 139229 73541
rect 139163 73476 139164 73540
rect 139228 73476 139229 73540
rect 139163 73475 139229 73476
rect 137794 71218 137826 71454
rect 138062 71218 138146 71454
rect 138382 71218 138414 71454
rect 137794 71134 138414 71218
rect 137794 70898 137826 71134
rect 138062 70898 138146 71134
rect 138382 70898 138414 71134
rect 137794 37454 138414 70898
rect 137794 37218 137826 37454
rect 138062 37218 138146 37454
rect 138382 37218 138414 37454
rect 137794 37134 138414 37218
rect 137794 36898 137826 37134
rect 138062 36898 138146 37134
rect 138382 36898 138414 37134
rect 137507 27028 137573 27029
rect 137507 26964 137508 27028
rect 137572 26964 137573 27028
rect 137507 26963 137573 26964
rect 133643 15876 133709 15877
rect 133643 15812 133644 15876
rect 133708 15812 133709 15876
rect 133643 15811 133709 15812
rect 137794 3454 138414 36898
rect 139166 25669 139226 73475
rect 139347 73404 139413 73405
rect 139347 73340 139348 73404
rect 139412 73340 139413 73404
rect 139347 73339 139413 73340
rect 140083 73404 140149 73405
rect 140083 73340 140084 73404
rect 140148 73340 140149 73404
rect 140083 73339 140149 73340
rect 139350 68373 139410 73339
rect 139347 68372 139413 68373
rect 139347 68308 139348 68372
rect 139412 68308 139413 68372
rect 139347 68307 139413 68308
rect 140086 54637 140146 73339
rect 140083 54636 140149 54637
rect 140083 54572 140084 54636
rect 140148 54572 140149 54636
rect 140083 54571 140149 54572
rect 140270 51917 140330 73611
rect 140451 73540 140517 73541
rect 140451 73476 140452 73540
rect 140516 73476 140517 73540
rect 140451 73475 140517 73476
rect 141187 73540 141253 73541
rect 141187 73476 141188 73540
rect 141252 73476 141253 73540
rect 141187 73475 141253 73476
rect 140267 51916 140333 51917
rect 140267 51852 140268 51916
rect 140332 51852 140333 51916
rect 140267 51851 140333 51852
rect 140454 36685 140514 73475
rect 140635 73404 140701 73405
rect 140635 73340 140636 73404
rect 140700 73340 140701 73404
rect 140635 73339 140701 73340
rect 140451 36684 140517 36685
rect 140451 36620 140452 36684
rect 140516 36620 140517 36684
rect 140451 36619 140517 36620
rect 139163 25668 139229 25669
rect 139163 25604 139164 25668
rect 139228 25604 139229 25668
rect 139163 25603 139229 25604
rect 140638 11933 140698 73339
rect 140635 11932 140701 11933
rect 140635 11868 140636 11932
rect 140700 11868 140701 11932
rect 140635 11867 140701 11868
rect 141190 3773 141250 73475
rect 141514 41174 142134 74063
rect 142843 72996 142909 72997
rect 142843 72932 142844 72996
rect 142908 72932 142909 72996
rect 142843 72931 142909 72932
rect 141514 40938 141546 41174
rect 141782 40938 141866 41174
rect 142102 40938 142134 41174
rect 141514 40854 142134 40938
rect 141514 40618 141546 40854
rect 141782 40618 141866 40854
rect 142102 40618 142134 40854
rect 141514 7174 142134 40618
rect 142846 19957 142906 72931
rect 143395 72860 143461 72861
rect 143395 72796 143396 72860
rect 143460 72796 143461 72860
rect 143395 72795 143461 72796
rect 144499 72860 144565 72861
rect 144499 72796 144500 72860
rect 144564 72796 144565 72860
rect 144499 72795 144565 72796
rect 145051 72860 145117 72861
rect 145051 72796 145052 72860
rect 145116 72796 145117 72860
rect 145051 72795 145117 72796
rect 143027 72724 143093 72725
rect 143027 72660 143028 72724
rect 143092 72660 143093 72724
rect 143027 72659 143093 72660
rect 143030 50421 143090 72659
rect 143211 72588 143277 72589
rect 143211 72524 143212 72588
rect 143276 72524 143277 72588
rect 143211 72523 143277 72524
rect 143027 50420 143093 50421
rect 143027 50356 143028 50420
rect 143092 50356 143093 50420
rect 143027 50355 143093 50356
rect 143214 49061 143274 72523
rect 143398 64293 143458 72795
rect 144315 72588 144381 72589
rect 144315 72524 144316 72588
rect 144380 72524 144381 72588
rect 144315 72523 144381 72524
rect 144131 72452 144197 72453
rect 144131 72388 144132 72452
rect 144196 72388 144197 72452
rect 144131 72387 144197 72388
rect 143395 64292 143461 64293
rect 143395 64228 143396 64292
rect 143460 64228 143461 64292
rect 143395 64227 143461 64228
rect 143211 49060 143277 49061
rect 143211 48996 143212 49060
rect 143276 48996 143277 49060
rect 143211 48995 143277 48996
rect 142843 19956 142909 19957
rect 142843 19892 142844 19956
rect 142908 19892 142909 19956
rect 142843 19891 142909 19892
rect 141514 6938 141546 7174
rect 141782 6938 141866 7174
rect 142102 6938 142134 7174
rect 141514 6854 142134 6938
rect 141514 6618 141546 6854
rect 141782 6618 141866 6854
rect 142102 6618 142134 6854
rect 141187 3772 141253 3773
rect 141187 3708 141188 3772
rect 141252 3708 141253 3772
rect 141187 3707 141253 3708
rect 132355 3364 132421 3365
rect 132355 3300 132356 3364
rect 132420 3300 132421 3364
rect 132355 3299 132421 3300
rect 129834 -7302 129866 -7066
rect 130102 -7302 130186 -7066
rect 130422 -7302 130454 -7066
rect 129834 -7386 130454 -7302
rect 129834 -7622 129866 -7386
rect 130102 -7622 130186 -7386
rect 130422 -7622 130454 -7386
rect 129834 -7654 130454 -7622
rect 137794 3218 137826 3454
rect 138062 3218 138146 3454
rect 138382 3218 138414 3454
rect 137794 3134 138414 3218
rect 137794 2898 137826 3134
rect 138062 2898 138146 3134
rect 138382 2898 138414 3134
rect 137794 -346 138414 2898
rect 137794 -582 137826 -346
rect 138062 -582 138146 -346
rect 138382 -582 138414 -346
rect 137794 -666 138414 -582
rect 137794 -902 137826 -666
rect 138062 -902 138146 -666
rect 138382 -902 138414 -666
rect 137794 -7654 138414 -902
rect 141514 -1306 142134 6618
rect 144134 3637 144194 72387
rect 144318 9077 144378 72523
rect 144315 9076 144381 9077
rect 144315 9012 144316 9076
rect 144380 9012 144381 9076
rect 144315 9011 144381 9012
rect 144131 3636 144197 3637
rect 144131 3572 144132 3636
rect 144196 3572 144197 3636
rect 144131 3571 144197 3572
rect 144502 3501 144562 72795
rect 144867 72724 144933 72725
rect 144867 72660 144868 72724
rect 144932 72660 144933 72724
rect 144867 72659 144933 72660
rect 144870 67013 144930 72659
rect 144867 67012 144933 67013
rect 144867 66948 144868 67012
rect 144932 66948 144933 67012
rect 144867 66947 144933 66948
rect 145054 58717 145114 72795
rect 145051 58716 145117 58717
rect 145051 58652 145052 58716
rect 145116 58652 145117 58716
rect 145051 58651 145117 58652
rect 145234 44894 145854 74063
rect 147446 73133 147506 75243
rect 160875 75172 160941 75173
rect 160875 75108 160876 75172
rect 160940 75108 160941 75172
rect 160875 75107 160941 75108
rect 158851 74900 158917 74901
rect 158851 74836 158852 74900
rect 158916 74836 158917 74900
rect 158851 74835 158917 74836
rect 155907 74764 155973 74765
rect 155907 74700 155908 74764
rect 155972 74700 155973 74764
rect 155907 74699 155973 74700
rect 147443 73132 147509 73133
rect 147443 73068 147444 73132
rect 147508 73068 147509 73132
rect 147443 73067 147509 73068
rect 147995 73132 148061 73133
rect 147995 73068 147996 73132
rect 148060 73068 148061 73132
rect 147995 73067 148061 73068
rect 147627 72996 147693 72997
rect 147627 72932 147628 72996
rect 147692 72932 147693 72996
rect 147627 72931 147693 72932
rect 146155 72724 146221 72725
rect 146155 72660 146156 72724
rect 146220 72660 146221 72724
rect 146155 72659 146221 72660
rect 147075 72724 147141 72725
rect 147075 72660 147076 72724
rect 147140 72660 147141 72724
rect 147075 72659 147141 72660
rect 145234 44658 145266 44894
rect 145502 44658 145586 44894
rect 145822 44658 145854 44894
rect 145234 44574 145854 44658
rect 145234 44338 145266 44574
rect 145502 44338 145586 44574
rect 145822 44338 145854 44574
rect 145234 10894 145854 44338
rect 145234 10658 145266 10894
rect 145502 10658 145586 10894
rect 145822 10658 145854 10894
rect 145234 10574 145854 10658
rect 145234 10338 145266 10574
rect 145502 10338 145586 10574
rect 145822 10338 145854 10574
rect 144499 3500 144565 3501
rect 144499 3436 144500 3500
rect 144564 3436 144565 3500
rect 144499 3435 144565 3436
rect 141514 -1542 141546 -1306
rect 141782 -1542 141866 -1306
rect 142102 -1542 142134 -1306
rect 141514 -1626 142134 -1542
rect 141514 -1862 141546 -1626
rect 141782 -1862 141866 -1626
rect 142102 -1862 142134 -1626
rect 141514 -7654 142134 -1862
rect 145234 -2266 145854 10338
rect 146158 8941 146218 72659
rect 146891 72180 146957 72181
rect 146891 72116 146892 72180
rect 146956 72116 146957 72180
rect 146891 72115 146957 72116
rect 146894 22813 146954 72115
rect 147078 47701 147138 72659
rect 147630 71909 147690 72931
rect 147627 71908 147693 71909
rect 147627 71844 147628 71908
rect 147692 71844 147693 71908
rect 147627 71843 147693 71844
rect 147443 71500 147509 71501
rect 147443 71436 147444 71500
rect 147508 71436 147509 71500
rect 147443 71435 147509 71436
rect 147259 71364 147325 71365
rect 147259 71300 147260 71364
rect 147324 71300 147325 71364
rect 147259 71299 147325 71300
rect 147075 47700 147141 47701
rect 147075 47636 147076 47700
rect 147140 47636 147141 47700
rect 147075 47635 147141 47636
rect 147262 46613 147322 71299
rect 147446 70410 147506 71435
rect 147446 70350 147874 70410
rect 147814 66877 147874 70350
rect 147811 66876 147877 66877
rect 147811 66812 147812 66876
rect 147876 66812 147877 66876
rect 147811 66811 147877 66812
rect 147259 46612 147325 46613
rect 147259 46548 147260 46612
rect 147324 46548 147325 46612
rect 147259 46547 147325 46548
rect 147998 44845 148058 73067
rect 148363 72860 148429 72861
rect 148363 72796 148364 72860
rect 148428 72796 148429 72860
rect 148363 72795 148429 72796
rect 148179 72588 148245 72589
rect 148179 72524 148180 72588
rect 148244 72524 148245 72588
rect 148179 72523 148245 72524
rect 147995 44844 148061 44845
rect 147995 44780 147996 44844
rect 148060 44780 148061 44844
rect 147995 44779 148061 44780
rect 148182 43485 148242 72523
rect 148179 43484 148245 43485
rect 148179 43420 148180 43484
rect 148244 43420 148245 43484
rect 148179 43419 148245 43420
rect 146891 22812 146957 22813
rect 146891 22748 146892 22812
rect 146956 22748 146957 22812
rect 146891 22747 146957 22748
rect 148366 21317 148426 72795
rect 148547 72724 148613 72725
rect 148547 72660 148548 72724
rect 148612 72660 148613 72724
rect 148547 72659 148613 72660
rect 148363 21316 148429 21317
rect 148363 21252 148364 21316
rect 148428 21252 148429 21316
rect 148363 21251 148429 21252
rect 148550 10301 148610 72659
rect 148954 48614 149574 74063
rect 151491 73948 151557 73949
rect 151491 73884 151492 73948
rect 151556 73884 151557 73948
rect 151491 73883 151557 73884
rect 150387 72860 150453 72861
rect 150387 72796 150388 72860
rect 150452 72796 150453 72860
rect 150387 72795 150453 72796
rect 150203 72724 150269 72725
rect 150203 72660 150204 72724
rect 150268 72660 150269 72724
rect 150203 72659 150269 72660
rect 148954 48378 148986 48614
rect 149222 48378 149306 48614
rect 149542 48378 149574 48614
rect 148954 48294 149574 48378
rect 148954 48058 148986 48294
rect 149222 48058 149306 48294
rect 149542 48058 149574 48294
rect 148954 14614 149574 48058
rect 150206 40765 150266 72659
rect 150390 69597 150450 72795
rect 151123 72588 151189 72589
rect 151123 72524 151124 72588
rect 151188 72524 151189 72588
rect 151123 72523 151189 72524
rect 150387 69596 150453 69597
rect 150387 69532 150388 69596
rect 150452 69532 150453 69596
rect 150387 69531 150453 69532
rect 151126 46477 151186 72523
rect 151307 72452 151373 72453
rect 151307 72388 151308 72452
rect 151372 72388 151373 72452
rect 151307 72387 151373 72388
rect 151123 46476 151189 46477
rect 151123 46412 151124 46476
rect 151188 46412 151189 46476
rect 151123 46411 151189 46412
rect 150203 40764 150269 40765
rect 150203 40700 150204 40764
rect 150268 40700 150269 40764
rect 150203 40699 150269 40700
rect 151310 39269 151370 72387
rect 151307 39268 151373 39269
rect 151307 39204 151308 39268
rect 151372 39204 151373 39268
rect 151307 39203 151373 39204
rect 151494 33829 151554 73883
rect 152227 72860 152293 72861
rect 152227 72796 152228 72860
rect 152292 72796 152293 72860
rect 152227 72795 152293 72796
rect 151675 72724 151741 72725
rect 151675 72660 151676 72724
rect 151740 72660 151741 72724
rect 151675 72659 151741 72660
rect 151491 33828 151557 33829
rect 151491 33764 151492 33828
rect 151556 33764 151557 33828
rect 151491 33763 151557 33764
rect 148954 14378 148986 14614
rect 149222 14378 149306 14614
rect 149542 14378 149574 14614
rect 148954 14294 149574 14378
rect 148954 14058 148986 14294
rect 149222 14058 149306 14294
rect 149542 14058 149574 14294
rect 148547 10300 148613 10301
rect 148547 10236 148548 10300
rect 148612 10236 148613 10300
rect 148547 10235 148613 10236
rect 146155 8940 146221 8941
rect 146155 8876 146156 8940
rect 146220 8876 146221 8940
rect 146155 8875 146221 8876
rect 145234 -2502 145266 -2266
rect 145502 -2502 145586 -2266
rect 145822 -2502 145854 -2266
rect 145234 -2586 145854 -2502
rect 145234 -2822 145266 -2586
rect 145502 -2822 145586 -2586
rect 145822 -2822 145854 -2586
rect 145234 -7654 145854 -2822
rect 148954 -3226 149574 14058
rect 151678 11797 151738 72659
rect 152230 37909 152290 72795
rect 152411 72724 152477 72725
rect 152411 72660 152412 72724
rect 152476 72660 152477 72724
rect 152411 72659 152477 72660
rect 152227 37908 152293 37909
rect 152227 37844 152228 37908
rect 152292 37844 152293 37908
rect 152227 37843 152293 37844
rect 152414 25533 152474 72659
rect 152674 52334 153294 74063
rect 153883 72860 153949 72861
rect 153883 72796 153884 72860
rect 153948 72796 153949 72860
rect 153883 72795 153949 72796
rect 155355 72860 155421 72861
rect 155355 72796 155356 72860
rect 155420 72796 155421 72860
rect 155355 72795 155421 72796
rect 152674 52098 152706 52334
rect 152942 52098 153026 52334
rect 153262 52098 153294 52334
rect 152674 52014 153294 52098
rect 152674 51778 152706 52014
rect 152942 51778 153026 52014
rect 153262 51778 153294 52014
rect 152411 25532 152477 25533
rect 152411 25468 152412 25532
rect 152476 25468 152477 25532
rect 152411 25467 152477 25468
rect 152674 18334 153294 51778
rect 153886 40629 153946 72795
rect 154251 72724 154317 72725
rect 154251 72660 154252 72724
rect 154316 72660 154317 72724
rect 154251 72659 154317 72660
rect 154067 72588 154133 72589
rect 154067 72524 154068 72588
rect 154132 72524 154133 72588
rect 154067 72523 154133 72524
rect 153883 40628 153949 40629
rect 153883 40564 153884 40628
rect 153948 40564 153949 40628
rect 153883 40563 153949 40564
rect 154070 36549 154130 72523
rect 154067 36548 154133 36549
rect 154067 36484 154068 36548
rect 154132 36484 154133 36548
rect 154067 36483 154133 36484
rect 154254 22677 154314 72659
rect 155171 72588 155237 72589
rect 155171 72524 155172 72588
rect 155236 72524 155237 72588
rect 155171 72523 155237 72524
rect 154435 72452 154501 72453
rect 154435 72388 154436 72452
rect 154500 72388 154501 72452
rect 154435 72387 154501 72388
rect 154251 22676 154317 22677
rect 154251 22612 154252 22676
rect 154316 22612 154317 22676
rect 154251 22611 154317 22612
rect 152674 18098 152706 18334
rect 152942 18098 153026 18334
rect 153262 18098 153294 18334
rect 152674 18014 153294 18098
rect 152674 17778 152706 18014
rect 152942 17778 153026 18014
rect 153262 17778 153294 18014
rect 151675 11796 151741 11797
rect 151675 11732 151676 11796
rect 151740 11732 151741 11796
rect 151675 11731 151741 11732
rect 148954 -3462 148986 -3226
rect 149222 -3462 149306 -3226
rect 149542 -3462 149574 -3226
rect 148954 -3546 149574 -3462
rect 148954 -3782 148986 -3546
rect 149222 -3782 149306 -3546
rect 149542 -3782 149574 -3546
rect 148954 -7654 149574 -3782
rect 152674 -4186 153294 17778
rect 154438 7581 154498 72387
rect 155174 59941 155234 72523
rect 155171 59940 155237 59941
rect 155171 59876 155172 59940
rect 155236 59876 155237 59940
rect 155171 59875 155237 59876
rect 155358 51781 155418 72795
rect 155723 72724 155789 72725
rect 155723 72660 155724 72724
rect 155788 72660 155789 72724
rect 155723 72659 155789 72660
rect 155539 72452 155605 72453
rect 155539 72388 155540 72452
rect 155604 72388 155605 72452
rect 155539 72387 155605 72388
rect 155355 51780 155421 51781
rect 155355 51716 155356 51780
rect 155420 51716 155421 51780
rect 155355 51715 155421 51716
rect 155542 35325 155602 72387
rect 155539 35324 155605 35325
rect 155539 35260 155540 35324
rect 155604 35260 155605 35324
rect 155539 35259 155605 35260
rect 155726 30973 155786 72659
rect 155910 71909 155970 74699
rect 157195 74628 157261 74629
rect 157195 74564 157196 74628
rect 157260 74564 157261 74628
rect 157195 74563 157261 74564
rect 155907 71908 155973 71909
rect 155907 71844 155908 71908
rect 155972 71844 155973 71908
rect 155907 71843 155973 71844
rect 156091 71908 156157 71909
rect 156091 71844 156092 71908
rect 156156 71844 156157 71908
rect 156091 71843 156157 71844
rect 156094 35189 156154 71843
rect 156394 56054 157014 74063
rect 157198 73949 157258 74563
rect 157195 73948 157261 73949
rect 157195 73884 157196 73948
rect 157260 73884 157261 73948
rect 157195 73883 157261 73884
rect 158854 73405 158914 74835
rect 158851 73404 158917 73405
rect 158851 73340 158852 73404
rect 158916 73340 158917 73404
rect 158851 73339 158917 73340
rect 157563 73132 157629 73133
rect 157563 73068 157564 73132
rect 157628 73068 157629 73132
rect 157563 73067 157629 73068
rect 157195 72588 157261 72589
rect 157195 72524 157196 72588
rect 157260 72524 157261 72588
rect 157195 72523 157261 72524
rect 156394 55818 156426 56054
rect 156662 55818 156746 56054
rect 156982 55818 157014 56054
rect 156394 55734 157014 55818
rect 156394 55498 156426 55734
rect 156662 55498 156746 55734
rect 156982 55498 157014 55734
rect 156091 35188 156157 35189
rect 156091 35124 156092 35188
rect 156156 35124 156157 35188
rect 156091 35123 156157 35124
rect 155723 30972 155789 30973
rect 155723 30908 155724 30972
rect 155788 30908 155789 30972
rect 155723 30907 155789 30908
rect 156394 22054 157014 55498
rect 156394 21818 156426 22054
rect 156662 21818 156746 22054
rect 156982 21818 157014 22054
rect 156394 21734 157014 21818
rect 156394 21498 156426 21734
rect 156662 21498 156746 21734
rect 156982 21498 157014 21734
rect 154435 7580 154501 7581
rect 154435 7516 154436 7580
rect 154500 7516 154501 7580
rect 154435 7515 154501 7516
rect 152674 -4422 152706 -4186
rect 152942 -4422 153026 -4186
rect 153262 -4422 153294 -4186
rect 152674 -4506 153294 -4422
rect 152674 -4742 152706 -4506
rect 152942 -4742 153026 -4506
rect 153262 -4742 153294 -4506
rect 152674 -7654 153294 -4742
rect 156394 -5146 157014 21498
rect 157198 3365 157258 72523
rect 157566 72181 157626 73067
rect 159035 72996 159101 72997
rect 159035 72932 159036 72996
rect 159100 72932 159101 72996
rect 159035 72931 159101 72932
rect 158299 72724 158365 72725
rect 158299 72660 158300 72724
rect 158364 72660 158365 72724
rect 158299 72659 158365 72660
rect 158667 72724 158733 72725
rect 158667 72660 158668 72724
rect 158732 72660 158733 72724
rect 158667 72659 158733 72660
rect 157931 72588 157997 72589
rect 157931 72524 157932 72588
rect 157996 72524 157997 72588
rect 157931 72523 157997 72524
rect 157747 72452 157813 72453
rect 157747 72388 157748 72452
rect 157812 72388 157813 72452
rect 157747 72387 157813 72388
rect 157563 72180 157629 72181
rect 157563 72116 157564 72180
rect 157628 72116 157629 72180
rect 157563 72115 157629 72116
rect 157750 57357 157810 72387
rect 157747 57356 157813 57357
rect 157747 57292 157748 57356
rect 157812 57292 157813 57356
rect 157747 57291 157813 57292
rect 157934 6221 157994 72523
rect 158302 6357 158362 72659
rect 158670 67149 158730 72659
rect 159038 72453 159098 72931
rect 159219 72724 159285 72725
rect 159219 72660 159220 72724
rect 159284 72660 159285 72724
rect 159219 72659 159285 72660
rect 159587 72724 159653 72725
rect 159587 72660 159588 72724
rect 159652 72660 159653 72724
rect 159587 72659 159653 72660
rect 159771 72724 159837 72725
rect 159771 72660 159772 72724
rect 159836 72660 159837 72724
rect 159771 72659 159837 72660
rect 159035 72452 159101 72453
rect 159035 72388 159036 72452
rect 159100 72388 159101 72452
rect 159035 72387 159101 72388
rect 158667 67148 158733 67149
rect 158667 67084 158668 67148
rect 158732 67084 158733 67148
rect 158667 67083 158733 67084
rect 159222 54501 159282 72659
rect 159403 72588 159469 72589
rect 159403 72524 159404 72588
rect 159468 72524 159469 72588
rect 159403 72523 159469 72524
rect 159219 54500 159285 54501
rect 159219 54436 159220 54500
rect 159284 54436 159285 54500
rect 159219 54435 159285 54436
rect 159406 26893 159466 72523
rect 159403 26892 159469 26893
rect 159403 26828 159404 26892
rect 159468 26828 159469 26892
rect 159403 26827 159469 26828
rect 159590 15877 159650 72659
rect 159587 15876 159653 15877
rect 159587 15812 159588 15876
rect 159652 15812 159653 15876
rect 159587 15811 159653 15812
rect 158299 6356 158365 6357
rect 158299 6292 158300 6356
rect 158364 6292 158365 6356
rect 158299 6291 158365 6292
rect 157931 6220 157997 6221
rect 157931 6156 157932 6220
rect 157996 6156 157997 6220
rect 157931 6155 157997 6156
rect 159774 4861 159834 72659
rect 160114 59774 160734 74063
rect 160878 72045 160938 75107
rect 161427 74900 161493 74901
rect 161427 74836 161428 74900
rect 161492 74836 161493 74900
rect 161427 74835 161493 74836
rect 161243 73268 161309 73269
rect 161243 73204 161244 73268
rect 161308 73204 161309 73268
rect 161243 73203 161309 73204
rect 161059 72588 161125 72589
rect 161059 72524 161060 72588
rect 161124 72524 161125 72588
rect 161059 72523 161125 72524
rect 160875 72044 160941 72045
rect 160875 71980 160876 72044
rect 160940 71980 160941 72044
rect 160875 71979 160941 71980
rect 160114 59538 160146 59774
rect 160382 59538 160466 59774
rect 160702 59538 160734 59774
rect 160114 59454 160734 59538
rect 160114 59218 160146 59454
rect 160382 59218 160466 59454
rect 160702 59218 160734 59454
rect 160114 25774 160734 59218
rect 161062 55861 161122 72523
rect 161059 55860 161125 55861
rect 161059 55796 161060 55860
rect 161124 55796 161125 55860
rect 161059 55795 161125 55796
rect 161246 50285 161306 73203
rect 161430 72317 161490 74835
rect 169342 74629 169402 75379
rect 169339 74628 169405 74629
rect 169339 74564 169340 74628
rect 169404 74564 169405 74628
rect 169339 74563 169405 74564
rect 161611 73540 161677 73541
rect 161611 73476 161612 73540
rect 161676 73476 161677 73540
rect 161611 73475 161677 73476
rect 161427 72316 161493 72317
rect 161427 72252 161428 72316
rect 161492 72252 161493 72316
rect 161427 72251 161493 72252
rect 161614 71365 161674 73475
rect 162163 73132 162229 73133
rect 162163 73068 162164 73132
rect 162228 73068 162229 73132
rect 162163 73067 162229 73068
rect 161611 71364 161677 71365
rect 161611 71300 161612 71364
rect 161676 71300 161677 71364
rect 161611 71299 161677 71300
rect 161243 50284 161309 50285
rect 161243 50220 161244 50284
rect 161308 50220 161309 50284
rect 161243 50219 161309 50220
rect 160114 25538 160146 25774
rect 160382 25538 160466 25774
rect 160702 25538 160734 25774
rect 160114 25454 160734 25538
rect 160114 25218 160146 25454
rect 160382 25218 160466 25454
rect 160702 25218 160734 25454
rect 159771 4860 159837 4861
rect 159771 4796 159772 4860
rect 159836 4796 159837 4860
rect 159771 4795 159837 4796
rect 157195 3364 157261 3365
rect 157195 3300 157196 3364
rect 157260 3300 157261 3364
rect 157195 3299 157261 3300
rect 156394 -5382 156426 -5146
rect 156662 -5382 156746 -5146
rect 156982 -5382 157014 -5146
rect 156394 -5466 157014 -5382
rect 156394 -5702 156426 -5466
rect 156662 -5702 156746 -5466
rect 156982 -5702 157014 -5466
rect 156394 -7654 157014 -5702
rect 160114 -6106 160734 25218
rect 162166 11661 162226 73067
rect 162531 72724 162597 72725
rect 162531 72660 162532 72724
rect 162596 72660 162597 72724
rect 162531 72659 162597 72660
rect 163451 72724 163517 72725
rect 163451 72660 163452 72724
rect 163516 72660 163517 72724
rect 163451 72659 163517 72660
rect 162347 72452 162413 72453
rect 162347 72388 162348 72452
rect 162412 72388 162413 72452
rect 162347 72387 162413 72388
rect 162350 57221 162410 72387
rect 162347 57220 162413 57221
rect 162347 57156 162348 57220
rect 162412 57156 162413 57220
rect 162347 57155 162413 57156
rect 162534 14517 162594 72659
rect 162715 72588 162781 72589
rect 162715 72524 162716 72588
rect 162780 72524 162781 72588
rect 162715 72523 162781 72524
rect 162718 65517 162778 72523
rect 163083 72452 163149 72453
rect 163083 72388 163084 72452
rect 163148 72388 163149 72452
rect 163083 72387 163149 72388
rect 163086 68237 163146 72387
rect 163083 68236 163149 68237
rect 163083 68172 163084 68236
rect 163148 68172 163149 68236
rect 163083 68171 163149 68172
rect 162715 65516 162781 65517
rect 162715 65452 162716 65516
rect 162780 65452 162781 65516
rect 162715 65451 162781 65452
rect 163454 42125 163514 72659
rect 163834 63494 164454 74063
rect 166211 73540 166277 73541
rect 166211 73476 166212 73540
rect 166276 73476 166277 73540
rect 166211 73475 166277 73476
rect 165291 72724 165357 72725
rect 165291 72660 165292 72724
rect 165356 72660 165357 72724
rect 165291 72659 165357 72660
rect 165107 72452 165173 72453
rect 165107 72388 165108 72452
rect 165172 72388 165173 72452
rect 165107 72387 165173 72388
rect 163834 63258 163866 63494
rect 164102 63258 164186 63494
rect 164422 63258 164454 63494
rect 163834 63174 164454 63258
rect 163834 62938 163866 63174
rect 164102 62938 164186 63174
rect 164422 62938 164454 63174
rect 163451 42124 163517 42125
rect 163451 42060 163452 42124
rect 163516 42060 163517 42124
rect 163451 42059 163517 42060
rect 163834 29494 164454 62938
rect 165110 48925 165170 72387
rect 165107 48924 165173 48925
rect 165107 48860 165108 48924
rect 165172 48860 165173 48924
rect 165107 48859 165173 48860
rect 165294 29613 165354 72659
rect 165475 72588 165541 72589
rect 165475 72524 165476 72588
rect 165540 72524 165541 72588
rect 165475 72523 165541 72524
rect 165291 29612 165357 29613
rect 165291 29548 165292 29612
rect 165356 29548 165357 29612
rect 165291 29547 165357 29548
rect 163834 29258 163866 29494
rect 164102 29258 164186 29494
rect 164422 29258 164454 29494
rect 163834 29174 164454 29258
rect 163834 28938 163866 29174
rect 164102 28938 164186 29174
rect 164422 28938 164454 29174
rect 162531 14516 162597 14517
rect 162531 14452 162532 14516
rect 162596 14452 162597 14516
rect 162531 14451 162597 14452
rect 162163 11660 162229 11661
rect 162163 11596 162164 11660
rect 162228 11596 162229 11660
rect 162163 11595 162229 11596
rect 160114 -6342 160146 -6106
rect 160382 -6342 160466 -6106
rect 160702 -6342 160734 -6106
rect 160114 -6426 160734 -6342
rect 160114 -6662 160146 -6426
rect 160382 -6662 160466 -6426
rect 160702 -6662 160734 -6426
rect 160114 -7654 160734 -6662
rect 163834 -7066 164454 28938
rect 165478 18733 165538 72523
rect 166214 71909 166274 73475
rect 166579 72588 166645 72589
rect 166579 72524 166580 72588
rect 166644 72524 166645 72588
rect 166579 72523 166645 72524
rect 166395 72180 166461 72181
rect 166395 72116 166396 72180
rect 166460 72116 166461 72180
rect 166395 72115 166461 72116
rect 166211 71908 166277 71909
rect 166211 71844 166212 71908
rect 166276 71844 166277 71908
rect 166211 71843 166277 71844
rect 166398 47565 166458 72115
rect 166395 47564 166461 47565
rect 166395 47500 166396 47564
rect 166460 47500 166461 47564
rect 166395 47499 166461 47500
rect 165475 18732 165541 18733
rect 165475 18668 165476 18732
rect 165540 18668 165541 18732
rect 165475 18667 165541 18668
rect 166582 18597 166642 72523
rect 166763 72452 166829 72453
rect 166763 72388 166764 72452
rect 166828 72388 166829 72452
rect 166763 72387 166829 72388
rect 166579 18596 166645 18597
rect 166579 18532 166580 18596
rect 166644 18532 166645 18596
rect 166579 18531 166645 18532
rect 166766 13021 166826 72387
rect 167499 72180 167565 72181
rect 167499 72116 167500 72180
rect 167564 72116 167565 72180
rect 167499 72115 167565 72116
rect 167502 46205 167562 72115
rect 171794 71454 172414 104898
rect 171794 71218 171826 71454
rect 172062 71218 172146 71454
rect 172382 71218 172414 71454
rect 171794 71134 172414 71218
rect 171794 70898 171826 71134
rect 172062 70898 172146 71134
rect 172382 70898 172414 71134
rect 167499 46204 167565 46205
rect 167499 46140 167500 46204
rect 167564 46140 167565 46204
rect 167499 46139 167565 46140
rect 171794 37454 172414 70898
rect 171794 37218 171826 37454
rect 172062 37218 172146 37454
rect 172382 37218 172414 37454
rect 171794 37134 172414 37218
rect 171794 36898 171826 37134
rect 172062 36898 172146 37134
rect 172382 36898 172414 37134
rect 166763 13020 166829 13021
rect 166763 12956 166764 13020
rect 166828 12956 166829 13020
rect 166763 12955 166829 12956
rect 163834 -7302 163866 -7066
rect 164102 -7302 164186 -7066
rect 164422 -7302 164454 -7066
rect 163834 -7386 164454 -7302
rect 163834 -7622 163866 -7386
rect 164102 -7622 164186 -7386
rect 164422 -7622 164454 -7386
rect 163834 -7654 164454 -7622
rect 171794 3454 172414 36898
rect 171794 3218 171826 3454
rect 172062 3218 172146 3454
rect 172382 3218 172414 3454
rect 171794 3134 172414 3218
rect 171794 2898 171826 3134
rect 172062 2898 172146 3134
rect 172382 2898 172414 3134
rect 171794 -346 172414 2898
rect 171794 -582 171826 -346
rect 172062 -582 172146 -346
rect 172382 -582 172414 -346
rect 171794 -666 172414 -582
rect 171794 -902 171826 -666
rect 172062 -902 172146 -666
rect 172382 -902 172414 -666
rect 171794 -7654 172414 -902
rect 175514 211174 176134 214340
rect 175514 210938 175546 211174
rect 175782 210938 175866 211174
rect 176102 210938 176134 211174
rect 175514 210854 176134 210938
rect 175514 210618 175546 210854
rect 175782 210618 175866 210854
rect 176102 210618 176134 210854
rect 175514 177174 176134 210618
rect 175514 176938 175546 177174
rect 175782 176938 175866 177174
rect 176102 176938 176134 177174
rect 175514 176854 176134 176938
rect 175514 176618 175546 176854
rect 175782 176618 175866 176854
rect 176102 176618 176134 176854
rect 175514 143174 176134 176618
rect 175514 142938 175546 143174
rect 175782 142938 175866 143174
rect 176102 142938 176134 143174
rect 175514 142854 176134 142938
rect 175514 142618 175546 142854
rect 175782 142618 175866 142854
rect 176102 142618 176134 142854
rect 175514 109174 176134 142618
rect 175514 108938 175546 109174
rect 175782 108938 175866 109174
rect 176102 108938 176134 109174
rect 175514 108854 176134 108938
rect 175514 108618 175546 108854
rect 175782 108618 175866 108854
rect 176102 108618 176134 108854
rect 175514 75174 176134 108618
rect 175514 74938 175546 75174
rect 175782 74938 175866 75174
rect 176102 74938 176134 75174
rect 175514 74854 176134 74938
rect 175514 74618 175546 74854
rect 175782 74618 175866 74854
rect 176102 74618 176134 74854
rect 175514 41174 176134 74618
rect 175514 40938 175546 41174
rect 175782 40938 175866 41174
rect 176102 40938 176134 41174
rect 175514 40854 176134 40938
rect 175514 40618 175546 40854
rect 175782 40618 175866 40854
rect 176102 40618 176134 40854
rect 175514 7174 176134 40618
rect 175514 6938 175546 7174
rect 175782 6938 175866 7174
rect 176102 6938 176134 7174
rect 175514 6854 176134 6938
rect 175514 6618 175546 6854
rect 175782 6618 175866 6854
rect 176102 6618 176134 6854
rect 175514 -1306 176134 6618
rect 175514 -1542 175546 -1306
rect 175782 -1542 175866 -1306
rect 176102 -1542 176134 -1306
rect 175514 -1626 176134 -1542
rect 175514 -1862 175546 -1626
rect 175782 -1862 175866 -1626
rect 176102 -1862 176134 -1626
rect 175514 -7654 176134 -1862
rect 179234 180894 179854 214340
rect 179234 180658 179266 180894
rect 179502 180658 179586 180894
rect 179822 180658 179854 180894
rect 179234 180574 179854 180658
rect 179234 180338 179266 180574
rect 179502 180338 179586 180574
rect 179822 180338 179854 180574
rect 179234 146894 179854 180338
rect 179234 146658 179266 146894
rect 179502 146658 179586 146894
rect 179822 146658 179854 146894
rect 179234 146574 179854 146658
rect 179234 146338 179266 146574
rect 179502 146338 179586 146574
rect 179822 146338 179854 146574
rect 179234 112894 179854 146338
rect 179234 112658 179266 112894
rect 179502 112658 179586 112894
rect 179822 112658 179854 112894
rect 179234 112574 179854 112658
rect 179234 112338 179266 112574
rect 179502 112338 179586 112574
rect 179822 112338 179854 112574
rect 179234 78894 179854 112338
rect 179234 78658 179266 78894
rect 179502 78658 179586 78894
rect 179822 78658 179854 78894
rect 179234 78574 179854 78658
rect 179234 78338 179266 78574
rect 179502 78338 179586 78574
rect 179822 78338 179854 78574
rect 179234 44894 179854 78338
rect 179234 44658 179266 44894
rect 179502 44658 179586 44894
rect 179822 44658 179854 44894
rect 179234 44574 179854 44658
rect 179234 44338 179266 44574
rect 179502 44338 179586 44574
rect 179822 44338 179854 44574
rect 179234 10894 179854 44338
rect 179234 10658 179266 10894
rect 179502 10658 179586 10894
rect 179822 10658 179854 10894
rect 179234 10574 179854 10658
rect 179234 10338 179266 10574
rect 179502 10338 179586 10574
rect 179822 10338 179854 10574
rect 179234 -2266 179854 10338
rect 179234 -2502 179266 -2266
rect 179502 -2502 179586 -2266
rect 179822 -2502 179854 -2266
rect 179234 -2586 179854 -2502
rect 179234 -2822 179266 -2586
rect 179502 -2822 179586 -2586
rect 179822 -2822 179854 -2586
rect 179234 -7654 179854 -2822
rect 182954 184614 183574 214340
rect 182954 184378 182986 184614
rect 183222 184378 183306 184614
rect 183542 184378 183574 184614
rect 182954 184294 183574 184378
rect 182954 184058 182986 184294
rect 183222 184058 183306 184294
rect 183542 184058 183574 184294
rect 182954 150614 183574 184058
rect 182954 150378 182986 150614
rect 183222 150378 183306 150614
rect 183542 150378 183574 150614
rect 182954 150294 183574 150378
rect 182954 150058 182986 150294
rect 183222 150058 183306 150294
rect 183542 150058 183574 150294
rect 182954 116614 183574 150058
rect 182954 116378 182986 116614
rect 183222 116378 183306 116614
rect 183542 116378 183574 116614
rect 182954 116294 183574 116378
rect 182954 116058 182986 116294
rect 183222 116058 183306 116294
rect 183542 116058 183574 116294
rect 182954 82614 183574 116058
rect 182954 82378 182986 82614
rect 183222 82378 183306 82614
rect 183542 82378 183574 82614
rect 182954 82294 183574 82378
rect 182954 82058 182986 82294
rect 183222 82058 183306 82294
rect 183542 82058 183574 82294
rect 182954 48614 183574 82058
rect 182954 48378 182986 48614
rect 183222 48378 183306 48614
rect 183542 48378 183574 48614
rect 182954 48294 183574 48378
rect 182954 48058 182986 48294
rect 183222 48058 183306 48294
rect 183542 48058 183574 48294
rect 182954 14614 183574 48058
rect 182954 14378 182986 14614
rect 183222 14378 183306 14614
rect 183542 14378 183574 14614
rect 182954 14294 183574 14378
rect 182954 14058 182986 14294
rect 183222 14058 183306 14294
rect 183542 14058 183574 14294
rect 182954 -3226 183574 14058
rect 182954 -3462 182986 -3226
rect 183222 -3462 183306 -3226
rect 183542 -3462 183574 -3226
rect 182954 -3546 183574 -3462
rect 182954 -3782 182986 -3546
rect 183222 -3782 183306 -3546
rect 183542 -3782 183574 -3546
rect 182954 -7654 183574 -3782
rect 186674 188334 187294 214340
rect 186674 188098 186706 188334
rect 186942 188098 187026 188334
rect 187262 188098 187294 188334
rect 186674 188014 187294 188098
rect 186674 187778 186706 188014
rect 186942 187778 187026 188014
rect 187262 187778 187294 188014
rect 186674 154334 187294 187778
rect 186674 154098 186706 154334
rect 186942 154098 187026 154334
rect 187262 154098 187294 154334
rect 186674 154014 187294 154098
rect 186674 153778 186706 154014
rect 186942 153778 187026 154014
rect 187262 153778 187294 154014
rect 186674 120334 187294 153778
rect 186674 120098 186706 120334
rect 186942 120098 187026 120334
rect 187262 120098 187294 120334
rect 186674 120014 187294 120098
rect 186674 119778 186706 120014
rect 186942 119778 187026 120014
rect 187262 119778 187294 120014
rect 186674 86334 187294 119778
rect 186674 86098 186706 86334
rect 186942 86098 187026 86334
rect 187262 86098 187294 86334
rect 186674 86014 187294 86098
rect 186674 85778 186706 86014
rect 186942 85778 187026 86014
rect 187262 85778 187294 86014
rect 186674 52334 187294 85778
rect 186674 52098 186706 52334
rect 186942 52098 187026 52334
rect 187262 52098 187294 52334
rect 186674 52014 187294 52098
rect 186674 51778 186706 52014
rect 186942 51778 187026 52014
rect 187262 51778 187294 52014
rect 186674 18334 187294 51778
rect 186674 18098 186706 18334
rect 186942 18098 187026 18334
rect 187262 18098 187294 18334
rect 186674 18014 187294 18098
rect 186674 17778 186706 18014
rect 186942 17778 187026 18014
rect 187262 17778 187294 18014
rect 186674 -4186 187294 17778
rect 186674 -4422 186706 -4186
rect 186942 -4422 187026 -4186
rect 187262 -4422 187294 -4186
rect 186674 -4506 187294 -4422
rect 186674 -4742 186706 -4506
rect 186942 -4742 187026 -4506
rect 187262 -4742 187294 -4506
rect 186674 -7654 187294 -4742
rect 190394 192054 191014 225498
rect 220674 222334 221294 255778
rect 224394 709638 225014 711590
rect 224394 709402 224426 709638
rect 224662 709402 224746 709638
rect 224982 709402 225014 709638
rect 224394 709318 225014 709402
rect 224394 709082 224426 709318
rect 224662 709082 224746 709318
rect 224982 709082 225014 709318
rect 224394 668054 225014 709082
rect 224394 667818 224426 668054
rect 224662 667818 224746 668054
rect 224982 667818 225014 668054
rect 224394 667734 225014 667818
rect 224394 667498 224426 667734
rect 224662 667498 224746 667734
rect 224982 667498 225014 667734
rect 224394 634054 225014 667498
rect 224394 633818 224426 634054
rect 224662 633818 224746 634054
rect 224982 633818 225014 634054
rect 224394 633734 225014 633818
rect 224394 633498 224426 633734
rect 224662 633498 224746 633734
rect 224982 633498 225014 633734
rect 224394 600054 225014 633498
rect 224394 599818 224426 600054
rect 224662 599818 224746 600054
rect 224982 599818 225014 600054
rect 224394 599734 225014 599818
rect 224394 599498 224426 599734
rect 224662 599498 224746 599734
rect 224982 599498 225014 599734
rect 224394 566054 225014 599498
rect 224394 565818 224426 566054
rect 224662 565818 224746 566054
rect 224982 565818 225014 566054
rect 224394 565734 225014 565818
rect 224394 565498 224426 565734
rect 224662 565498 224746 565734
rect 224982 565498 225014 565734
rect 224394 532054 225014 565498
rect 224394 531818 224426 532054
rect 224662 531818 224746 532054
rect 224982 531818 225014 532054
rect 224394 531734 225014 531818
rect 224394 531498 224426 531734
rect 224662 531498 224746 531734
rect 224982 531498 225014 531734
rect 224394 498054 225014 531498
rect 224394 497818 224426 498054
rect 224662 497818 224746 498054
rect 224982 497818 225014 498054
rect 224394 497734 225014 497818
rect 224394 497498 224426 497734
rect 224662 497498 224746 497734
rect 224982 497498 225014 497734
rect 224394 464054 225014 497498
rect 224394 463818 224426 464054
rect 224662 463818 224746 464054
rect 224982 463818 225014 464054
rect 224394 463734 225014 463818
rect 224394 463498 224426 463734
rect 224662 463498 224746 463734
rect 224982 463498 225014 463734
rect 224394 430054 225014 463498
rect 224394 429818 224426 430054
rect 224662 429818 224746 430054
rect 224982 429818 225014 430054
rect 224394 429734 225014 429818
rect 224394 429498 224426 429734
rect 224662 429498 224746 429734
rect 224982 429498 225014 429734
rect 224394 396054 225014 429498
rect 224394 395818 224426 396054
rect 224662 395818 224746 396054
rect 224982 395818 225014 396054
rect 224394 395734 225014 395818
rect 224394 395498 224426 395734
rect 224662 395498 224746 395734
rect 224982 395498 225014 395734
rect 224394 362054 225014 395498
rect 224394 361818 224426 362054
rect 224662 361818 224746 362054
rect 224982 361818 225014 362054
rect 224394 361734 225014 361818
rect 224394 361498 224426 361734
rect 224662 361498 224746 361734
rect 224982 361498 225014 361734
rect 224394 328054 225014 361498
rect 224394 327818 224426 328054
rect 224662 327818 224746 328054
rect 224982 327818 225014 328054
rect 224394 327734 225014 327818
rect 224394 327498 224426 327734
rect 224662 327498 224746 327734
rect 224982 327498 225014 327734
rect 224394 294054 225014 327498
rect 224394 293818 224426 294054
rect 224662 293818 224746 294054
rect 224982 293818 225014 294054
rect 224394 293734 225014 293818
rect 224394 293498 224426 293734
rect 224662 293498 224746 293734
rect 224982 293498 225014 293734
rect 224394 260054 225014 293498
rect 224394 259818 224426 260054
rect 224662 259818 224746 260054
rect 224982 259818 225014 260054
rect 224394 259734 225014 259818
rect 224394 259498 224426 259734
rect 224662 259498 224746 259734
rect 224982 259498 225014 259734
rect 224394 225991 225014 259498
rect 224394 225755 224426 225991
rect 224662 225755 224746 225991
rect 224982 225755 225014 225991
rect 224394 225660 225014 225755
rect 228114 710598 228734 711590
rect 228114 710362 228146 710598
rect 228382 710362 228466 710598
rect 228702 710362 228734 710598
rect 228114 710278 228734 710362
rect 228114 710042 228146 710278
rect 228382 710042 228466 710278
rect 228702 710042 228734 710278
rect 228114 671774 228734 710042
rect 228114 671538 228146 671774
rect 228382 671538 228466 671774
rect 228702 671538 228734 671774
rect 228114 671454 228734 671538
rect 228114 671218 228146 671454
rect 228382 671218 228466 671454
rect 228702 671218 228734 671454
rect 228114 637774 228734 671218
rect 228114 637538 228146 637774
rect 228382 637538 228466 637774
rect 228702 637538 228734 637774
rect 228114 637454 228734 637538
rect 228114 637218 228146 637454
rect 228382 637218 228466 637454
rect 228702 637218 228734 637454
rect 228114 603774 228734 637218
rect 228114 603538 228146 603774
rect 228382 603538 228466 603774
rect 228702 603538 228734 603774
rect 228114 603454 228734 603538
rect 228114 603218 228146 603454
rect 228382 603218 228466 603454
rect 228702 603218 228734 603454
rect 228114 569774 228734 603218
rect 228114 569538 228146 569774
rect 228382 569538 228466 569774
rect 228702 569538 228734 569774
rect 228114 569454 228734 569538
rect 228114 569218 228146 569454
rect 228382 569218 228466 569454
rect 228702 569218 228734 569454
rect 228114 535774 228734 569218
rect 228114 535538 228146 535774
rect 228382 535538 228466 535774
rect 228702 535538 228734 535774
rect 228114 535454 228734 535538
rect 228114 535218 228146 535454
rect 228382 535218 228466 535454
rect 228702 535218 228734 535454
rect 228114 501774 228734 535218
rect 228114 501538 228146 501774
rect 228382 501538 228466 501774
rect 228702 501538 228734 501774
rect 228114 501454 228734 501538
rect 228114 501218 228146 501454
rect 228382 501218 228466 501454
rect 228702 501218 228734 501454
rect 228114 467774 228734 501218
rect 228114 467538 228146 467774
rect 228382 467538 228466 467774
rect 228702 467538 228734 467774
rect 228114 467454 228734 467538
rect 228114 467218 228146 467454
rect 228382 467218 228466 467454
rect 228702 467218 228734 467454
rect 228114 433774 228734 467218
rect 228114 433538 228146 433774
rect 228382 433538 228466 433774
rect 228702 433538 228734 433774
rect 228114 433454 228734 433538
rect 228114 433218 228146 433454
rect 228382 433218 228466 433454
rect 228702 433218 228734 433454
rect 228114 399774 228734 433218
rect 228114 399538 228146 399774
rect 228382 399538 228466 399774
rect 228702 399538 228734 399774
rect 228114 399454 228734 399538
rect 228114 399218 228146 399454
rect 228382 399218 228466 399454
rect 228702 399218 228734 399454
rect 228114 365774 228734 399218
rect 228114 365538 228146 365774
rect 228382 365538 228466 365774
rect 228702 365538 228734 365774
rect 228114 365454 228734 365538
rect 228114 365218 228146 365454
rect 228382 365218 228466 365454
rect 228702 365218 228734 365454
rect 228114 331774 228734 365218
rect 228114 331538 228146 331774
rect 228382 331538 228466 331774
rect 228702 331538 228734 331774
rect 228114 331454 228734 331538
rect 228114 331218 228146 331454
rect 228382 331218 228466 331454
rect 228702 331218 228734 331454
rect 228114 297774 228734 331218
rect 228114 297538 228146 297774
rect 228382 297538 228466 297774
rect 228702 297538 228734 297774
rect 228114 297454 228734 297538
rect 228114 297218 228146 297454
rect 228382 297218 228466 297454
rect 228702 297218 228734 297454
rect 228114 263774 228734 297218
rect 228114 263538 228146 263774
rect 228382 263538 228466 263774
rect 228702 263538 228734 263774
rect 228114 263454 228734 263538
rect 228114 263218 228146 263454
rect 228382 263218 228466 263454
rect 228702 263218 228734 263454
rect 228114 229774 228734 263218
rect 228114 229538 228146 229774
rect 228382 229538 228466 229774
rect 228702 229538 228734 229774
rect 228114 229454 228734 229538
rect 228114 229218 228146 229454
rect 228382 229218 228466 229454
rect 228702 229218 228734 229454
rect 228114 225660 228734 229218
rect 231834 711558 232454 711590
rect 231834 711322 231866 711558
rect 232102 711322 232186 711558
rect 232422 711322 232454 711558
rect 231834 711238 232454 711322
rect 231834 711002 231866 711238
rect 232102 711002 232186 711238
rect 232422 711002 232454 711238
rect 231834 675494 232454 711002
rect 231834 675258 231866 675494
rect 232102 675258 232186 675494
rect 232422 675258 232454 675494
rect 231834 675174 232454 675258
rect 231834 674938 231866 675174
rect 232102 674938 232186 675174
rect 232422 674938 232454 675174
rect 231834 641494 232454 674938
rect 231834 641258 231866 641494
rect 232102 641258 232186 641494
rect 232422 641258 232454 641494
rect 231834 641174 232454 641258
rect 231834 640938 231866 641174
rect 232102 640938 232186 641174
rect 232422 640938 232454 641174
rect 231834 607494 232454 640938
rect 231834 607258 231866 607494
rect 232102 607258 232186 607494
rect 232422 607258 232454 607494
rect 231834 607174 232454 607258
rect 231834 606938 231866 607174
rect 232102 606938 232186 607174
rect 232422 606938 232454 607174
rect 231834 573494 232454 606938
rect 231834 573258 231866 573494
rect 232102 573258 232186 573494
rect 232422 573258 232454 573494
rect 231834 573174 232454 573258
rect 231834 572938 231866 573174
rect 232102 572938 232186 573174
rect 232422 572938 232454 573174
rect 231834 539494 232454 572938
rect 231834 539258 231866 539494
rect 232102 539258 232186 539494
rect 232422 539258 232454 539494
rect 231834 539174 232454 539258
rect 231834 538938 231866 539174
rect 232102 538938 232186 539174
rect 232422 538938 232454 539174
rect 231834 505494 232454 538938
rect 231834 505258 231866 505494
rect 232102 505258 232186 505494
rect 232422 505258 232454 505494
rect 231834 505174 232454 505258
rect 231834 504938 231866 505174
rect 232102 504938 232186 505174
rect 232422 504938 232454 505174
rect 231834 471494 232454 504938
rect 231834 471258 231866 471494
rect 232102 471258 232186 471494
rect 232422 471258 232454 471494
rect 231834 471174 232454 471258
rect 231834 470938 231866 471174
rect 232102 470938 232186 471174
rect 232422 470938 232454 471174
rect 231834 437494 232454 470938
rect 231834 437258 231866 437494
rect 232102 437258 232186 437494
rect 232422 437258 232454 437494
rect 231834 437174 232454 437258
rect 231834 436938 231866 437174
rect 232102 436938 232186 437174
rect 232422 436938 232454 437174
rect 231834 403494 232454 436938
rect 231834 403258 231866 403494
rect 232102 403258 232186 403494
rect 232422 403258 232454 403494
rect 231834 403174 232454 403258
rect 231834 402938 231866 403174
rect 232102 402938 232186 403174
rect 232422 402938 232454 403174
rect 231834 369494 232454 402938
rect 231834 369258 231866 369494
rect 232102 369258 232186 369494
rect 232422 369258 232454 369494
rect 231834 369174 232454 369258
rect 231834 368938 231866 369174
rect 232102 368938 232186 369174
rect 232422 368938 232454 369174
rect 231834 335494 232454 368938
rect 231834 335258 231866 335494
rect 232102 335258 232186 335494
rect 232422 335258 232454 335494
rect 231834 335174 232454 335258
rect 231834 334938 231866 335174
rect 232102 334938 232186 335174
rect 232422 334938 232454 335174
rect 231834 301494 232454 334938
rect 231834 301258 231866 301494
rect 232102 301258 232186 301494
rect 232422 301258 232454 301494
rect 231834 301174 232454 301258
rect 231834 300938 231866 301174
rect 232102 300938 232186 301174
rect 232422 300938 232454 301174
rect 231834 267494 232454 300938
rect 231834 267258 231866 267494
rect 232102 267258 232186 267494
rect 232422 267258 232454 267494
rect 231834 267174 232454 267258
rect 231834 266938 231866 267174
rect 232102 266938 232186 267174
rect 232422 266938 232454 267174
rect 231834 233494 232454 266938
rect 231834 233258 231866 233494
rect 232102 233258 232186 233494
rect 232422 233258 232454 233494
rect 231834 233174 232454 233258
rect 231834 232938 231866 233174
rect 232102 232938 232186 233174
rect 232422 232938 232454 233174
rect 231834 225660 232454 232938
rect 239794 704838 240414 711590
rect 239794 704602 239826 704838
rect 240062 704602 240146 704838
rect 240382 704602 240414 704838
rect 239794 704518 240414 704602
rect 239794 704282 239826 704518
rect 240062 704282 240146 704518
rect 240382 704282 240414 704518
rect 239794 683454 240414 704282
rect 239794 683218 239826 683454
rect 240062 683218 240146 683454
rect 240382 683218 240414 683454
rect 239794 683134 240414 683218
rect 239794 682898 239826 683134
rect 240062 682898 240146 683134
rect 240382 682898 240414 683134
rect 239794 649454 240414 682898
rect 239794 649218 239826 649454
rect 240062 649218 240146 649454
rect 240382 649218 240414 649454
rect 239794 649134 240414 649218
rect 239794 648898 239826 649134
rect 240062 648898 240146 649134
rect 240382 648898 240414 649134
rect 239794 615454 240414 648898
rect 239794 615218 239826 615454
rect 240062 615218 240146 615454
rect 240382 615218 240414 615454
rect 239794 615134 240414 615218
rect 239794 614898 239826 615134
rect 240062 614898 240146 615134
rect 240382 614898 240414 615134
rect 239794 581454 240414 614898
rect 239794 581218 239826 581454
rect 240062 581218 240146 581454
rect 240382 581218 240414 581454
rect 239794 581134 240414 581218
rect 239794 580898 239826 581134
rect 240062 580898 240146 581134
rect 240382 580898 240414 581134
rect 239794 547454 240414 580898
rect 239794 547218 239826 547454
rect 240062 547218 240146 547454
rect 240382 547218 240414 547454
rect 239794 547134 240414 547218
rect 239794 546898 239826 547134
rect 240062 546898 240146 547134
rect 240382 546898 240414 547134
rect 239794 513454 240414 546898
rect 239794 513218 239826 513454
rect 240062 513218 240146 513454
rect 240382 513218 240414 513454
rect 239794 513134 240414 513218
rect 239794 512898 239826 513134
rect 240062 512898 240146 513134
rect 240382 512898 240414 513134
rect 239794 479454 240414 512898
rect 239794 479218 239826 479454
rect 240062 479218 240146 479454
rect 240382 479218 240414 479454
rect 239794 479134 240414 479218
rect 239794 478898 239826 479134
rect 240062 478898 240146 479134
rect 240382 478898 240414 479134
rect 239794 445454 240414 478898
rect 239794 445218 239826 445454
rect 240062 445218 240146 445454
rect 240382 445218 240414 445454
rect 239794 445134 240414 445218
rect 239794 444898 239826 445134
rect 240062 444898 240146 445134
rect 240382 444898 240414 445134
rect 239794 411454 240414 444898
rect 239794 411218 239826 411454
rect 240062 411218 240146 411454
rect 240382 411218 240414 411454
rect 239794 411134 240414 411218
rect 239794 410898 239826 411134
rect 240062 410898 240146 411134
rect 240382 410898 240414 411134
rect 239794 377454 240414 410898
rect 239794 377218 239826 377454
rect 240062 377218 240146 377454
rect 240382 377218 240414 377454
rect 239794 377134 240414 377218
rect 239794 376898 239826 377134
rect 240062 376898 240146 377134
rect 240382 376898 240414 377134
rect 239794 343454 240414 376898
rect 239794 343218 239826 343454
rect 240062 343218 240146 343454
rect 240382 343218 240414 343454
rect 239794 343134 240414 343218
rect 239794 342898 239826 343134
rect 240062 342898 240146 343134
rect 240382 342898 240414 343134
rect 239794 309454 240414 342898
rect 239794 309218 239826 309454
rect 240062 309218 240146 309454
rect 240382 309218 240414 309454
rect 239794 309134 240414 309218
rect 239794 308898 239826 309134
rect 240062 308898 240146 309134
rect 240382 308898 240414 309134
rect 239794 275454 240414 308898
rect 239794 275218 239826 275454
rect 240062 275218 240146 275454
rect 240382 275218 240414 275454
rect 239794 275134 240414 275218
rect 239794 274898 239826 275134
rect 240062 274898 240146 275134
rect 240382 274898 240414 275134
rect 239794 241454 240414 274898
rect 239794 241218 239826 241454
rect 240062 241218 240146 241454
rect 240382 241218 240414 241454
rect 239794 241134 240414 241218
rect 239794 240898 239826 241134
rect 240062 240898 240146 241134
rect 240382 240898 240414 241134
rect 239794 225660 240414 240898
rect 243514 705798 244134 711590
rect 243514 705562 243546 705798
rect 243782 705562 243866 705798
rect 244102 705562 244134 705798
rect 243514 705478 244134 705562
rect 243514 705242 243546 705478
rect 243782 705242 243866 705478
rect 244102 705242 244134 705478
rect 243514 687174 244134 705242
rect 243514 686938 243546 687174
rect 243782 686938 243866 687174
rect 244102 686938 244134 687174
rect 243514 686854 244134 686938
rect 243514 686618 243546 686854
rect 243782 686618 243866 686854
rect 244102 686618 244134 686854
rect 243514 653174 244134 686618
rect 243514 652938 243546 653174
rect 243782 652938 243866 653174
rect 244102 652938 244134 653174
rect 243514 652854 244134 652938
rect 243514 652618 243546 652854
rect 243782 652618 243866 652854
rect 244102 652618 244134 652854
rect 243514 619174 244134 652618
rect 243514 618938 243546 619174
rect 243782 618938 243866 619174
rect 244102 618938 244134 619174
rect 243514 618854 244134 618938
rect 243514 618618 243546 618854
rect 243782 618618 243866 618854
rect 244102 618618 244134 618854
rect 243514 585174 244134 618618
rect 243514 584938 243546 585174
rect 243782 584938 243866 585174
rect 244102 584938 244134 585174
rect 243514 584854 244134 584938
rect 243514 584618 243546 584854
rect 243782 584618 243866 584854
rect 244102 584618 244134 584854
rect 243514 551174 244134 584618
rect 243514 550938 243546 551174
rect 243782 550938 243866 551174
rect 244102 550938 244134 551174
rect 243514 550854 244134 550938
rect 243514 550618 243546 550854
rect 243782 550618 243866 550854
rect 244102 550618 244134 550854
rect 243514 517174 244134 550618
rect 243514 516938 243546 517174
rect 243782 516938 243866 517174
rect 244102 516938 244134 517174
rect 243514 516854 244134 516938
rect 243514 516618 243546 516854
rect 243782 516618 243866 516854
rect 244102 516618 244134 516854
rect 243514 483174 244134 516618
rect 243514 482938 243546 483174
rect 243782 482938 243866 483174
rect 244102 482938 244134 483174
rect 243514 482854 244134 482938
rect 243514 482618 243546 482854
rect 243782 482618 243866 482854
rect 244102 482618 244134 482854
rect 243514 449174 244134 482618
rect 243514 448938 243546 449174
rect 243782 448938 243866 449174
rect 244102 448938 244134 449174
rect 243514 448854 244134 448938
rect 243514 448618 243546 448854
rect 243782 448618 243866 448854
rect 244102 448618 244134 448854
rect 243514 415174 244134 448618
rect 243514 414938 243546 415174
rect 243782 414938 243866 415174
rect 244102 414938 244134 415174
rect 243514 414854 244134 414938
rect 243514 414618 243546 414854
rect 243782 414618 243866 414854
rect 244102 414618 244134 414854
rect 243514 381174 244134 414618
rect 243514 380938 243546 381174
rect 243782 380938 243866 381174
rect 244102 380938 244134 381174
rect 243514 380854 244134 380938
rect 243514 380618 243546 380854
rect 243782 380618 243866 380854
rect 244102 380618 244134 380854
rect 243514 347174 244134 380618
rect 243514 346938 243546 347174
rect 243782 346938 243866 347174
rect 244102 346938 244134 347174
rect 243514 346854 244134 346938
rect 243514 346618 243546 346854
rect 243782 346618 243866 346854
rect 244102 346618 244134 346854
rect 243514 313174 244134 346618
rect 243514 312938 243546 313174
rect 243782 312938 243866 313174
rect 244102 312938 244134 313174
rect 243514 312854 244134 312938
rect 243514 312618 243546 312854
rect 243782 312618 243866 312854
rect 244102 312618 244134 312854
rect 243514 279174 244134 312618
rect 243514 278938 243546 279174
rect 243782 278938 243866 279174
rect 244102 278938 244134 279174
rect 243514 278854 244134 278938
rect 243514 278618 243546 278854
rect 243782 278618 243866 278854
rect 244102 278618 244134 278854
rect 243514 245174 244134 278618
rect 243514 244938 243546 245174
rect 243782 244938 243866 245174
rect 244102 244938 244134 245174
rect 243514 244854 244134 244938
rect 243514 244618 243546 244854
rect 243782 244618 243866 244854
rect 244102 244618 244134 244854
rect 243514 225660 244134 244618
rect 247234 706758 247854 711590
rect 247234 706522 247266 706758
rect 247502 706522 247586 706758
rect 247822 706522 247854 706758
rect 247234 706438 247854 706522
rect 247234 706202 247266 706438
rect 247502 706202 247586 706438
rect 247822 706202 247854 706438
rect 247234 690894 247854 706202
rect 247234 690658 247266 690894
rect 247502 690658 247586 690894
rect 247822 690658 247854 690894
rect 247234 690574 247854 690658
rect 247234 690338 247266 690574
rect 247502 690338 247586 690574
rect 247822 690338 247854 690574
rect 247234 656894 247854 690338
rect 247234 656658 247266 656894
rect 247502 656658 247586 656894
rect 247822 656658 247854 656894
rect 247234 656574 247854 656658
rect 247234 656338 247266 656574
rect 247502 656338 247586 656574
rect 247822 656338 247854 656574
rect 247234 622894 247854 656338
rect 247234 622658 247266 622894
rect 247502 622658 247586 622894
rect 247822 622658 247854 622894
rect 247234 622574 247854 622658
rect 247234 622338 247266 622574
rect 247502 622338 247586 622574
rect 247822 622338 247854 622574
rect 247234 588894 247854 622338
rect 247234 588658 247266 588894
rect 247502 588658 247586 588894
rect 247822 588658 247854 588894
rect 247234 588574 247854 588658
rect 247234 588338 247266 588574
rect 247502 588338 247586 588574
rect 247822 588338 247854 588574
rect 247234 554894 247854 588338
rect 247234 554658 247266 554894
rect 247502 554658 247586 554894
rect 247822 554658 247854 554894
rect 247234 554574 247854 554658
rect 247234 554338 247266 554574
rect 247502 554338 247586 554574
rect 247822 554338 247854 554574
rect 247234 520894 247854 554338
rect 247234 520658 247266 520894
rect 247502 520658 247586 520894
rect 247822 520658 247854 520894
rect 247234 520574 247854 520658
rect 247234 520338 247266 520574
rect 247502 520338 247586 520574
rect 247822 520338 247854 520574
rect 247234 486894 247854 520338
rect 247234 486658 247266 486894
rect 247502 486658 247586 486894
rect 247822 486658 247854 486894
rect 247234 486574 247854 486658
rect 247234 486338 247266 486574
rect 247502 486338 247586 486574
rect 247822 486338 247854 486574
rect 247234 452894 247854 486338
rect 247234 452658 247266 452894
rect 247502 452658 247586 452894
rect 247822 452658 247854 452894
rect 247234 452574 247854 452658
rect 247234 452338 247266 452574
rect 247502 452338 247586 452574
rect 247822 452338 247854 452574
rect 247234 418894 247854 452338
rect 247234 418658 247266 418894
rect 247502 418658 247586 418894
rect 247822 418658 247854 418894
rect 247234 418574 247854 418658
rect 247234 418338 247266 418574
rect 247502 418338 247586 418574
rect 247822 418338 247854 418574
rect 247234 384894 247854 418338
rect 247234 384658 247266 384894
rect 247502 384658 247586 384894
rect 247822 384658 247854 384894
rect 247234 384574 247854 384658
rect 247234 384338 247266 384574
rect 247502 384338 247586 384574
rect 247822 384338 247854 384574
rect 247234 350894 247854 384338
rect 247234 350658 247266 350894
rect 247502 350658 247586 350894
rect 247822 350658 247854 350894
rect 247234 350574 247854 350658
rect 247234 350338 247266 350574
rect 247502 350338 247586 350574
rect 247822 350338 247854 350574
rect 247234 316894 247854 350338
rect 247234 316658 247266 316894
rect 247502 316658 247586 316894
rect 247822 316658 247854 316894
rect 247234 316574 247854 316658
rect 247234 316338 247266 316574
rect 247502 316338 247586 316574
rect 247822 316338 247854 316574
rect 247234 282894 247854 316338
rect 247234 282658 247266 282894
rect 247502 282658 247586 282894
rect 247822 282658 247854 282894
rect 247234 282574 247854 282658
rect 247234 282338 247266 282574
rect 247502 282338 247586 282574
rect 247822 282338 247854 282574
rect 247234 248894 247854 282338
rect 247234 248658 247266 248894
rect 247502 248658 247586 248894
rect 247822 248658 247854 248894
rect 247234 248574 247854 248658
rect 247234 248338 247266 248574
rect 247502 248338 247586 248574
rect 247822 248338 247854 248574
rect 247234 225660 247854 248338
rect 250954 707718 251574 711590
rect 250954 707482 250986 707718
rect 251222 707482 251306 707718
rect 251542 707482 251574 707718
rect 250954 707398 251574 707482
rect 250954 707162 250986 707398
rect 251222 707162 251306 707398
rect 251542 707162 251574 707398
rect 250954 694614 251574 707162
rect 250954 694378 250986 694614
rect 251222 694378 251306 694614
rect 251542 694378 251574 694614
rect 250954 694294 251574 694378
rect 250954 694058 250986 694294
rect 251222 694058 251306 694294
rect 251542 694058 251574 694294
rect 250954 660614 251574 694058
rect 250954 660378 250986 660614
rect 251222 660378 251306 660614
rect 251542 660378 251574 660614
rect 250954 660294 251574 660378
rect 250954 660058 250986 660294
rect 251222 660058 251306 660294
rect 251542 660058 251574 660294
rect 250954 626614 251574 660058
rect 250954 626378 250986 626614
rect 251222 626378 251306 626614
rect 251542 626378 251574 626614
rect 250954 626294 251574 626378
rect 250954 626058 250986 626294
rect 251222 626058 251306 626294
rect 251542 626058 251574 626294
rect 250954 592614 251574 626058
rect 250954 592378 250986 592614
rect 251222 592378 251306 592614
rect 251542 592378 251574 592614
rect 250954 592294 251574 592378
rect 250954 592058 250986 592294
rect 251222 592058 251306 592294
rect 251542 592058 251574 592294
rect 250954 558614 251574 592058
rect 250954 558378 250986 558614
rect 251222 558378 251306 558614
rect 251542 558378 251574 558614
rect 250954 558294 251574 558378
rect 250954 558058 250986 558294
rect 251222 558058 251306 558294
rect 251542 558058 251574 558294
rect 250954 524614 251574 558058
rect 250954 524378 250986 524614
rect 251222 524378 251306 524614
rect 251542 524378 251574 524614
rect 250954 524294 251574 524378
rect 250954 524058 250986 524294
rect 251222 524058 251306 524294
rect 251542 524058 251574 524294
rect 250954 490614 251574 524058
rect 250954 490378 250986 490614
rect 251222 490378 251306 490614
rect 251542 490378 251574 490614
rect 250954 490294 251574 490378
rect 250954 490058 250986 490294
rect 251222 490058 251306 490294
rect 251542 490058 251574 490294
rect 250954 456614 251574 490058
rect 250954 456378 250986 456614
rect 251222 456378 251306 456614
rect 251542 456378 251574 456614
rect 250954 456294 251574 456378
rect 250954 456058 250986 456294
rect 251222 456058 251306 456294
rect 251542 456058 251574 456294
rect 250954 422614 251574 456058
rect 250954 422378 250986 422614
rect 251222 422378 251306 422614
rect 251542 422378 251574 422614
rect 250954 422294 251574 422378
rect 250954 422058 250986 422294
rect 251222 422058 251306 422294
rect 251542 422058 251574 422294
rect 250954 388614 251574 422058
rect 250954 388378 250986 388614
rect 251222 388378 251306 388614
rect 251542 388378 251574 388614
rect 250954 388294 251574 388378
rect 250954 388058 250986 388294
rect 251222 388058 251306 388294
rect 251542 388058 251574 388294
rect 250954 354614 251574 388058
rect 250954 354378 250986 354614
rect 251222 354378 251306 354614
rect 251542 354378 251574 354614
rect 250954 354294 251574 354378
rect 250954 354058 250986 354294
rect 251222 354058 251306 354294
rect 251542 354058 251574 354294
rect 250954 320614 251574 354058
rect 250954 320378 250986 320614
rect 251222 320378 251306 320614
rect 251542 320378 251574 320614
rect 250954 320294 251574 320378
rect 250954 320058 250986 320294
rect 251222 320058 251306 320294
rect 251542 320058 251574 320294
rect 250954 286614 251574 320058
rect 250954 286378 250986 286614
rect 251222 286378 251306 286614
rect 251542 286378 251574 286614
rect 250954 286294 251574 286378
rect 250954 286058 250986 286294
rect 251222 286058 251306 286294
rect 251542 286058 251574 286294
rect 250954 252614 251574 286058
rect 250954 252378 250986 252614
rect 251222 252378 251306 252614
rect 251542 252378 251574 252614
rect 250954 252294 251574 252378
rect 250954 252058 250986 252294
rect 251222 252058 251306 252294
rect 251542 252058 251574 252294
rect 220674 222098 220706 222334
rect 220942 222098 221026 222334
rect 221262 222098 221294 222334
rect 220674 222014 221294 222098
rect 220674 221778 220706 222014
rect 220942 221778 221026 222014
rect 221262 221778 221294 222014
rect 190394 191818 190426 192054
rect 190662 191818 190746 192054
rect 190982 191818 191014 192054
rect 190394 191734 191014 191818
rect 190394 191498 190426 191734
rect 190662 191498 190746 191734
rect 190982 191498 191014 191734
rect 190394 158054 191014 191498
rect 190394 157818 190426 158054
rect 190662 157818 190746 158054
rect 190982 157818 191014 158054
rect 190394 157734 191014 157818
rect 190394 157498 190426 157734
rect 190662 157498 190746 157734
rect 190982 157498 191014 157734
rect 190394 124054 191014 157498
rect 190394 123818 190426 124054
rect 190662 123818 190746 124054
rect 190982 123818 191014 124054
rect 190394 123734 191014 123818
rect 190394 123498 190426 123734
rect 190662 123498 190746 123734
rect 190982 123498 191014 123734
rect 190394 90054 191014 123498
rect 190394 89818 190426 90054
rect 190662 89818 190746 90054
rect 190982 89818 191014 90054
rect 190394 89734 191014 89818
rect 190394 89498 190426 89734
rect 190662 89498 190746 89734
rect 190982 89498 191014 89734
rect 190394 56054 191014 89498
rect 190394 55818 190426 56054
rect 190662 55818 190746 56054
rect 190982 55818 191014 56054
rect 190394 55734 191014 55818
rect 190394 55498 190426 55734
rect 190662 55498 190746 55734
rect 190982 55498 191014 55734
rect 190394 22054 191014 55498
rect 190394 21818 190426 22054
rect 190662 21818 190746 22054
rect 190982 21818 191014 22054
rect 190394 21734 191014 21818
rect 190394 21498 190426 21734
rect 190662 21498 190746 21734
rect 190982 21498 191014 21734
rect 190394 -5146 191014 21498
rect 190394 -5382 190426 -5146
rect 190662 -5382 190746 -5146
rect 190982 -5382 191014 -5146
rect 190394 -5466 191014 -5382
rect 190394 -5702 190426 -5466
rect 190662 -5702 190746 -5466
rect 190982 -5702 191014 -5466
rect 190394 -7654 191014 -5702
rect 194114 195774 194734 214340
rect 194114 195538 194146 195774
rect 194382 195538 194466 195774
rect 194702 195538 194734 195774
rect 194114 195454 194734 195538
rect 194114 195218 194146 195454
rect 194382 195218 194466 195454
rect 194702 195218 194734 195454
rect 194114 161774 194734 195218
rect 194114 161538 194146 161774
rect 194382 161538 194466 161774
rect 194702 161538 194734 161774
rect 194114 161454 194734 161538
rect 194114 161218 194146 161454
rect 194382 161218 194466 161454
rect 194702 161218 194734 161454
rect 194114 127774 194734 161218
rect 194114 127538 194146 127774
rect 194382 127538 194466 127774
rect 194702 127538 194734 127774
rect 194114 127454 194734 127538
rect 194114 127218 194146 127454
rect 194382 127218 194466 127454
rect 194702 127218 194734 127454
rect 194114 93774 194734 127218
rect 194114 93538 194146 93774
rect 194382 93538 194466 93774
rect 194702 93538 194734 93774
rect 194114 93454 194734 93538
rect 194114 93218 194146 93454
rect 194382 93218 194466 93454
rect 194702 93218 194734 93454
rect 194114 59774 194734 93218
rect 194114 59538 194146 59774
rect 194382 59538 194466 59774
rect 194702 59538 194734 59774
rect 194114 59454 194734 59538
rect 194114 59218 194146 59454
rect 194382 59218 194466 59454
rect 194702 59218 194734 59454
rect 194114 25774 194734 59218
rect 194114 25538 194146 25774
rect 194382 25538 194466 25774
rect 194702 25538 194734 25774
rect 194114 25454 194734 25538
rect 194114 25218 194146 25454
rect 194382 25218 194466 25454
rect 194702 25218 194734 25454
rect 194114 -6106 194734 25218
rect 194114 -6342 194146 -6106
rect 194382 -6342 194466 -6106
rect 194702 -6342 194734 -6106
rect 194114 -6426 194734 -6342
rect 194114 -6662 194146 -6426
rect 194382 -6662 194466 -6426
rect 194702 -6662 194734 -6426
rect 194114 -7654 194734 -6662
rect 197834 199494 198454 214340
rect 197834 199258 197866 199494
rect 198102 199258 198186 199494
rect 198422 199258 198454 199494
rect 197834 199174 198454 199258
rect 197834 198938 197866 199174
rect 198102 198938 198186 199174
rect 198422 198938 198454 199174
rect 197834 165494 198454 198938
rect 197834 165258 197866 165494
rect 198102 165258 198186 165494
rect 198422 165258 198454 165494
rect 197834 165174 198454 165258
rect 197834 164938 197866 165174
rect 198102 164938 198186 165174
rect 198422 164938 198454 165174
rect 197834 131494 198454 164938
rect 197834 131258 197866 131494
rect 198102 131258 198186 131494
rect 198422 131258 198454 131494
rect 197834 131174 198454 131258
rect 197834 130938 197866 131174
rect 198102 130938 198186 131174
rect 198422 130938 198454 131174
rect 197834 97494 198454 130938
rect 197834 97258 197866 97494
rect 198102 97258 198186 97494
rect 198422 97258 198454 97494
rect 197834 97174 198454 97258
rect 197834 96938 197866 97174
rect 198102 96938 198186 97174
rect 198422 96938 198454 97174
rect 197834 63494 198454 96938
rect 197834 63258 197866 63494
rect 198102 63258 198186 63494
rect 198422 63258 198454 63494
rect 197834 63174 198454 63258
rect 197834 62938 197866 63174
rect 198102 62938 198186 63174
rect 198422 62938 198454 63174
rect 197834 29494 198454 62938
rect 197834 29258 197866 29494
rect 198102 29258 198186 29494
rect 198422 29258 198454 29494
rect 197834 29174 198454 29258
rect 197834 28938 197866 29174
rect 198102 28938 198186 29174
rect 198422 28938 198454 29174
rect 197834 -7066 198454 28938
rect 197834 -7302 197866 -7066
rect 198102 -7302 198186 -7066
rect 198422 -7302 198454 -7066
rect 197834 -7386 198454 -7302
rect 197834 -7622 197866 -7386
rect 198102 -7622 198186 -7386
rect 198422 -7622 198454 -7386
rect 197834 -7654 198454 -7622
rect 205794 207454 206414 214340
rect 205794 207218 205826 207454
rect 206062 207218 206146 207454
rect 206382 207218 206414 207454
rect 205794 207134 206414 207218
rect 205794 206898 205826 207134
rect 206062 206898 206146 207134
rect 206382 206898 206414 207134
rect 205794 173454 206414 206898
rect 205794 173218 205826 173454
rect 206062 173218 206146 173454
rect 206382 173218 206414 173454
rect 205794 173134 206414 173218
rect 205794 172898 205826 173134
rect 206062 172898 206146 173134
rect 206382 172898 206414 173134
rect 205794 139454 206414 172898
rect 205794 139218 205826 139454
rect 206062 139218 206146 139454
rect 206382 139218 206414 139454
rect 205794 139134 206414 139218
rect 205794 138898 205826 139134
rect 206062 138898 206146 139134
rect 206382 138898 206414 139134
rect 205794 105454 206414 138898
rect 205794 105218 205826 105454
rect 206062 105218 206146 105454
rect 206382 105218 206414 105454
rect 205794 105134 206414 105218
rect 205794 104898 205826 105134
rect 206062 104898 206146 105134
rect 206382 104898 206414 105134
rect 205794 71454 206414 104898
rect 205794 71218 205826 71454
rect 206062 71218 206146 71454
rect 206382 71218 206414 71454
rect 205794 71134 206414 71218
rect 205794 70898 205826 71134
rect 206062 70898 206146 71134
rect 206382 70898 206414 71134
rect 205794 37454 206414 70898
rect 205794 37218 205826 37454
rect 206062 37218 206146 37454
rect 206382 37218 206414 37454
rect 205794 37134 206414 37218
rect 205794 36898 205826 37134
rect 206062 36898 206146 37134
rect 206382 36898 206414 37134
rect 205794 3454 206414 36898
rect 205794 3218 205826 3454
rect 206062 3218 206146 3454
rect 206382 3218 206414 3454
rect 205794 3134 206414 3218
rect 205794 2898 205826 3134
rect 206062 2898 206146 3134
rect 206382 2898 206414 3134
rect 205794 -346 206414 2898
rect 205794 -582 205826 -346
rect 206062 -582 206146 -346
rect 206382 -582 206414 -346
rect 205794 -666 206414 -582
rect 205794 -902 205826 -666
rect 206062 -902 206146 -666
rect 206382 -902 206414 -666
rect 205794 -7654 206414 -902
rect 209514 211174 210134 214340
rect 209514 210938 209546 211174
rect 209782 210938 209866 211174
rect 210102 210938 210134 211174
rect 209514 210854 210134 210938
rect 209514 210618 209546 210854
rect 209782 210618 209866 210854
rect 210102 210618 210134 210854
rect 209514 177174 210134 210618
rect 209514 176938 209546 177174
rect 209782 176938 209866 177174
rect 210102 176938 210134 177174
rect 209514 176854 210134 176938
rect 209514 176618 209546 176854
rect 209782 176618 209866 176854
rect 210102 176618 210134 176854
rect 209514 143174 210134 176618
rect 209514 142938 209546 143174
rect 209782 142938 209866 143174
rect 210102 142938 210134 143174
rect 209514 142854 210134 142938
rect 209514 142618 209546 142854
rect 209782 142618 209866 142854
rect 210102 142618 210134 142854
rect 209514 109174 210134 142618
rect 209514 108938 209546 109174
rect 209782 108938 209866 109174
rect 210102 108938 210134 109174
rect 209514 108854 210134 108938
rect 209514 108618 209546 108854
rect 209782 108618 209866 108854
rect 210102 108618 210134 108854
rect 209514 75174 210134 108618
rect 209514 74938 209546 75174
rect 209782 74938 209866 75174
rect 210102 74938 210134 75174
rect 209514 74854 210134 74938
rect 209514 74618 209546 74854
rect 209782 74618 209866 74854
rect 210102 74618 210134 74854
rect 209514 41174 210134 74618
rect 209514 40938 209546 41174
rect 209782 40938 209866 41174
rect 210102 40938 210134 41174
rect 209514 40854 210134 40938
rect 209514 40618 209546 40854
rect 209782 40618 209866 40854
rect 210102 40618 210134 40854
rect 209514 7174 210134 40618
rect 209514 6938 209546 7174
rect 209782 6938 209866 7174
rect 210102 6938 210134 7174
rect 209514 6854 210134 6938
rect 209514 6618 209546 6854
rect 209782 6618 209866 6854
rect 210102 6618 210134 6854
rect 209514 -1306 210134 6618
rect 209514 -1542 209546 -1306
rect 209782 -1542 209866 -1306
rect 210102 -1542 210134 -1306
rect 209514 -1626 210134 -1542
rect 209514 -1862 209546 -1626
rect 209782 -1862 209866 -1626
rect 210102 -1862 210134 -1626
rect 209514 -7654 210134 -1862
rect 213234 180894 213854 214340
rect 213234 180658 213266 180894
rect 213502 180658 213586 180894
rect 213822 180658 213854 180894
rect 213234 180574 213854 180658
rect 213234 180338 213266 180574
rect 213502 180338 213586 180574
rect 213822 180338 213854 180574
rect 213234 146894 213854 180338
rect 213234 146658 213266 146894
rect 213502 146658 213586 146894
rect 213822 146658 213854 146894
rect 213234 146574 213854 146658
rect 213234 146338 213266 146574
rect 213502 146338 213586 146574
rect 213822 146338 213854 146574
rect 213234 112894 213854 146338
rect 213234 112658 213266 112894
rect 213502 112658 213586 112894
rect 213822 112658 213854 112894
rect 213234 112574 213854 112658
rect 213234 112338 213266 112574
rect 213502 112338 213586 112574
rect 213822 112338 213854 112574
rect 213234 78894 213854 112338
rect 213234 78658 213266 78894
rect 213502 78658 213586 78894
rect 213822 78658 213854 78894
rect 213234 78574 213854 78658
rect 213234 78338 213266 78574
rect 213502 78338 213586 78574
rect 213822 78338 213854 78574
rect 213234 44894 213854 78338
rect 213234 44658 213266 44894
rect 213502 44658 213586 44894
rect 213822 44658 213854 44894
rect 213234 44574 213854 44658
rect 213234 44338 213266 44574
rect 213502 44338 213586 44574
rect 213822 44338 213854 44574
rect 213234 10894 213854 44338
rect 213234 10658 213266 10894
rect 213502 10658 213586 10894
rect 213822 10658 213854 10894
rect 213234 10574 213854 10658
rect 213234 10338 213266 10574
rect 213502 10338 213586 10574
rect 213822 10338 213854 10574
rect 213234 -2266 213854 10338
rect 213234 -2502 213266 -2266
rect 213502 -2502 213586 -2266
rect 213822 -2502 213854 -2266
rect 213234 -2586 213854 -2502
rect 213234 -2822 213266 -2586
rect 213502 -2822 213586 -2586
rect 213822 -2822 213854 -2586
rect 213234 -7654 213854 -2822
rect 216954 184614 217574 214340
rect 216954 184378 216986 184614
rect 217222 184378 217306 184614
rect 217542 184378 217574 184614
rect 216954 184294 217574 184378
rect 216954 184058 216986 184294
rect 217222 184058 217306 184294
rect 217542 184058 217574 184294
rect 216954 150614 217574 184058
rect 216954 150378 216986 150614
rect 217222 150378 217306 150614
rect 217542 150378 217574 150614
rect 216954 150294 217574 150378
rect 216954 150058 216986 150294
rect 217222 150058 217306 150294
rect 217542 150058 217574 150294
rect 216954 116614 217574 150058
rect 216954 116378 216986 116614
rect 217222 116378 217306 116614
rect 217542 116378 217574 116614
rect 216954 116294 217574 116378
rect 216954 116058 216986 116294
rect 217222 116058 217306 116294
rect 217542 116058 217574 116294
rect 216954 82614 217574 116058
rect 216954 82378 216986 82614
rect 217222 82378 217306 82614
rect 217542 82378 217574 82614
rect 216954 82294 217574 82378
rect 216954 82058 216986 82294
rect 217222 82058 217306 82294
rect 217542 82058 217574 82294
rect 216954 48614 217574 82058
rect 216954 48378 216986 48614
rect 217222 48378 217306 48614
rect 217542 48378 217574 48614
rect 216954 48294 217574 48378
rect 216954 48058 216986 48294
rect 217222 48058 217306 48294
rect 217542 48058 217574 48294
rect 216954 14614 217574 48058
rect 216954 14378 216986 14614
rect 217222 14378 217306 14614
rect 217542 14378 217574 14614
rect 216954 14294 217574 14378
rect 216954 14058 216986 14294
rect 217222 14058 217306 14294
rect 217542 14058 217574 14294
rect 216954 -3226 217574 14058
rect 216954 -3462 216986 -3226
rect 217222 -3462 217306 -3226
rect 217542 -3462 217574 -3226
rect 216954 -3546 217574 -3462
rect 216954 -3782 216986 -3546
rect 217222 -3782 217306 -3546
rect 217542 -3782 217574 -3546
rect 216954 -7654 217574 -3782
rect 220674 188334 221294 221778
rect 250954 218614 251574 252058
rect 254674 708678 255294 711590
rect 254674 708442 254706 708678
rect 254942 708442 255026 708678
rect 255262 708442 255294 708678
rect 254674 708358 255294 708442
rect 254674 708122 254706 708358
rect 254942 708122 255026 708358
rect 255262 708122 255294 708358
rect 254674 698334 255294 708122
rect 254674 698098 254706 698334
rect 254942 698098 255026 698334
rect 255262 698098 255294 698334
rect 254674 698014 255294 698098
rect 254674 697778 254706 698014
rect 254942 697778 255026 698014
rect 255262 697778 255294 698014
rect 254674 664334 255294 697778
rect 254674 664098 254706 664334
rect 254942 664098 255026 664334
rect 255262 664098 255294 664334
rect 254674 664014 255294 664098
rect 254674 663778 254706 664014
rect 254942 663778 255026 664014
rect 255262 663778 255294 664014
rect 254674 630334 255294 663778
rect 254674 630098 254706 630334
rect 254942 630098 255026 630334
rect 255262 630098 255294 630334
rect 254674 630014 255294 630098
rect 254674 629778 254706 630014
rect 254942 629778 255026 630014
rect 255262 629778 255294 630014
rect 254674 596334 255294 629778
rect 254674 596098 254706 596334
rect 254942 596098 255026 596334
rect 255262 596098 255294 596334
rect 254674 596014 255294 596098
rect 254674 595778 254706 596014
rect 254942 595778 255026 596014
rect 255262 595778 255294 596014
rect 254674 562334 255294 595778
rect 254674 562098 254706 562334
rect 254942 562098 255026 562334
rect 255262 562098 255294 562334
rect 254674 562014 255294 562098
rect 254674 561778 254706 562014
rect 254942 561778 255026 562014
rect 255262 561778 255294 562014
rect 254674 528334 255294 561778
rect 254674 528098 254706 528334
rect 254942 528098 255026 528334
rect 255262 528098 255294 528334
rect 254674 528014 255294 528098
rect 254674 527778 254706 528014
rect 254942 527778 255026 528014
rect 255262 527778 255294 528014
rect 254674 494334 255294 527778
rect 254674 494098 254706 494334
rect 254942 494098 255026 494334
rect 255262 494098 255294 494334
rect 254674 494014 255294 494098
rect 254674 493778 254706 494014
rect 254942 493778 255026 494014
rect 255262 493778 255294 494014
rect 254674 460334 255294 493778
rect 254674 460098 254706 460334
rect 254942 460098 255026 460334
rect 255262 460098 255294 460334
rect 254674 460014 255294 460098
rect 254674 459778 254706 460014
rect 254942 459778 255026 460014
rect 255262 459778 255294 460014
rect 254674 426334 255294 459778
rect 254674 426098 254706 426334
rect 254942 426098 255026 426334
rect 255262 426098 255294 426334
rect 254674 426014 255294 426098
rect 254674 425778 254706 426014
rect 254942 425778 255026 426014
rect 255262 425778 255294 426014
rect 254674 392334 255294 425778
rect 254674 392098 254706 392334
rect 254942 392098 255026 392334
rect 255262 392098 255294 392334
rect 254674 392014 255294 392098
rect 254674 391778 254706 392014
rect 254942 391778 255026 392014
rect 255262 391778 255294 392014
rect 254674 358334 255294 391778
rect 254674 358098 254706 358334
rect 254942 358098 255026 358334
rect 255262 358098 255294 358334
rect 254674 358014 255294 358098
rect 254674 357778 254706 358014
rect 254942 357778 255026 358014
rect 255262 357778 255294 358014
rect 254674 324334 255294 357778
rect 254674 324098 254706 324334
rect 254942 324098 255026 324334
rect 255262 324098 255294 324334
rect 254674 324014 255294 324098
rect 254674 323778 254706 324014
rect 254942 323778 255026 324014
rect 255262 323778 255294 324014
rect 254674 290334 255294 323778
rect 254674 290098 254706 290334
rect 254942 290098 255026 290334
rect 255262 290098 255294 290334
rect 254674 290014 255294 290098
rect 254674 289778 254706 290014
rect 254942 289778 255026 290014
rect 255262 289778 255294 290014
rect 254674 256334 255294 289778
rect 254674 256098 254706 256334
rect 254942 256098 255026 256334
rect 255262 256098 255294 256334
rect 254674 256014 255294 256098
rect 254674 255778 254706 256014
rect 254942 255778 255026 256014
rect 255262 255778 255294 256014
rect 254674 225660 255294 255778
rect 258394 709638 259014 711590
rect 258394 709402 258426 709638
rect 258662 709402 258746 709638
rect 258982 709402 259014 709638
rect 258394 709318 259014 709402
rect 258394 709082 258426 709318
rect 258662 709082 258746 709318
rect 258982 709082 259014 709318
rect 258394 668054 259014 709082
rect 258394 667818 258426 668054
rect 258662 667818 258746 668054
rect 258982 667818 259014 668054
rect 258394 667734 259014 667818
rect 258394 667498 258426 667734
rect 258662 667498 258746 667734
rect 258982 667498 259014 667734
rect 258394 634054 259014 667498
rect 258394 633818 258426 634054
rect 258662 633818 258746 634054
rect 258982 633818 259014 634054
rect 258394 633734 259014 633818
rect 258394 633498 258426 633734
rect 258662 633498 258746 633734
rect 258982 633498 259014 633734
rect 258394 600054 259014 633498
rect 258394 599818 258426 600054
rect 258662 599818 258746 600054
rect 258982 599818 259014 600054
rect 258394 599734 259014 599818
rect 258394 599498 258426 599734
rect 258662 599498 258746 599734
rect 258982 599498 259014 599734
rect 258394 566054 259014 599498
rect 258394 565818 258426 566054
rect 258662 565818 258746 566054
rect 258982 565818 259014 566054
rect 258394 565734 259014 565818
rect 258394 565498 258426 565734
rect 258662 565498 258746 565734
rect 258982 565498 259014 565734
rect 258394 532054 259014 565498
rect 258394 531818 258426 532054
rect 258662 531818 258746 532054
rect 258982 531818 259014 532054
rect 258394 531734 259014 531818
rect 258394 531498 258426 531734
rect 258662 531498 258746 531734
rect 258982 531498 259014 531734
rect 258394 498054 259014 531498
rect 258394 497818 258426 498054
rect 258662 497818 258746 498054
rect 258982 497818 259014 498054
rect 258394 497734 259014 497818
rect 258394 497498 258426 497734
rect 258662 497498 258746 497734
rect 258982 497498 259014 497734
rect 258394 464054 259014 497498
rect 258394 463818 258426 464054
rect 258662 463818 258746 464054
rect 258982 463818 259014 464054
rect 258394 463734 259014 463818
rect 258394 463498 258426 463734
rect 258662 463498 258746 463734
rect 258982 463498 259014 463734
rect 258394 430054 259014 463498
rect 258394 429818 258426 430054
rect 258662 429818 258746 430054
rect 258982 429818 259014 430054
rect 258394 429734 259014 429818
rect 258394 429498 258426 429734
rect 258662 429498 258746 429734
rect 258982 429498 259014 429734
rect 258394 396054 259014 429498
rect 258394 395818 258426 396054
rect 258662 395818 258746 396054
rect 258982 395818 259014 396054
rect 258394 395734 259014 395818
rect 258394 395498 258426 395734
rect 258662 395498 258746 395734
rect 258982 395498 259014 395734
rect 258394 362054 259014 395498
rect 258394 361818 258426 362054
rect 258662 361818 258746 362054
rect 258982 361818 259014 362054
rect 258394 361734 259014 361818
rect 258394 361498 258426 361734
rect 258662 361498 258746 361734
rect 258982 361498 259014 361734
rect 258394 328054 259014 361498
rect 258394 327818 258426 328054
rect 258662 327818 258746 328054
rect 258982 327818 259014 328054
rect 258394 327734 259014 327818
rect 258394 327498 258426 327734
rect 258662 327498 258746 327734
rect 258982 327498 259014 327734
rect 258394 294054 259014 327498
rect 258394 293818 258426 294054
rect 258662 293818 258746 294054
rect 258982 293818 259014 294054
rect 258394 293734 259014 293818
rect 258394 293498 258426 293734
rect 258662 293498 258746 293734
rect 258982 293498 259014 293734
rect 258394 260054 259014 293498
rect 258394 259818 258426 260054
rect 258662 259818 258746 260054
rect 258982 259818 259014 260054
rect 258394 259734 259014 259818
rect 258394 259498 258426 259734
rect 258662 259498 258746 259734
rect 258982 259498 259014 259734
rect 258394 225991 259014 259498
rect 258394 225755 258426 225991
rect 258662 225755 258746 225991
rect 258982 225755 259014 225991
rect 258394 225660 259014 225755
rect 262114 710598 262734 711590
rect 262114 710362 262146 710598
rect 262382 710362 262466 710598
rect 262702 710362 262734 710598
rect 262114 710278 262734 710362
rect 262114 710042 262146 710278
rect 262382 710042 262466 710278
rect 262702 710042 262734 710278
rect 262114 671774 262734 710042
rect 262114 671538 262146 671774
rect 262382 671538 262466 671774
rect 262702 671538 262734 671774
rect 262114 671454 262734 671538
rect 262114 671218 262146 671454
rect 262382 671218 262466 671454
rect 262702 671218 262734 671454
rect 262114 637774 262734 671218
rect 262114 637538 262146 637774
rect 262382 637538 262466 637774
rect 262702 637538 262734 637774
rect 262114 637454 262734 637538
rect 262114 637218 262146 637454
rect 262382 637218 262466 637454
rect 262702 637218 262734 637454
rect 262114 603774 262734 637218
rect 262114 603538 262146 603774
rect 262382 603538 262466 603774
rect 262702 603538 262734 603774
rect 262114 603454 262734 603538
rect 262114 603218 262146 603454
rect 262382 603218 262466 603454
rect 262702 603218 262734 603454
rect 262114 569774 262734 603218
rect 262114 569538 262146 569774
rect 262382 569538 262466 569774
rect 262702 569538 262734 569774
rect 262114 569454 262734 569538
rect 262114 569218 262146 569454
rect 262382 569218 262466 569454
rect 262702 569218 262734 569454
rect 262114 535774 262734 569218
rect 262114 535538 262146 535774
rect 262382 535538 262466 535774
rect 262702 535538 262734 535774
rect 262114 535454 262734 535538
rect 262114 535218 262146 535454
rect 262382 535218 262466 535454
rect 262702 535218 262734 535454
rect 262114 501774 262734 535218
rect 262114 501538 262146 501774
rect 262382 501538 262466 501774
rect 262702 501538 262734 501774
rect 262114 501454 262734 501538
rect 262114 501218 262146 501454
rect 262382 501218 262466 501454
rect 262702 501218 262734 501454
rect 262114 467774 262734 501218
rect 262114 467538 262146 467774
rect 262382 467538 262466 467774
rect 262702 467538 262734 467774
rect 262114 467454 262734 467538
rect 262114 467218 262146 467454
rect 262382 467218 262466 467454
rect 262702 467218 262734 467454
rect 262114 433774 262734 467218
rect 262114 433538 262146 433774
rect 262382 433538 262466 433774
rect 262702 433538 262734 433774
rect 262114 433454 262734 433538
rect 262114 433218 262146 433454
rect 262382 433218 262466 433454
rect 262702 433218 262734 433454
rect 262114 399774 262734 433218
rect 262114 399538 262146 399774
rect 262382 399538 262466 399774
rect 262702 399538 262734 399774
rect 262114 399454 262734 399538
rect 262114 399218 262146 399454
rect 262382 399218 262466 399454
rect 262702 399218 262734 399454
rect 262114 365774 262734 399218
rect 262114 365538 262146 365774
rect 262382 365538 262466 365774
rect 262702 365538 262734 365774
rect 262114 365454 262734 365538
rect 262114 365218 262146 365454
rect 262382 365218 262466 365454
rect 262702 365218 262734 365454
rect 262114 331774 262734 365218
rect 262114 331538 262146 331774
rect 262382 331538 262466 331774
rect 262702 331538 262734 331774
rect 262114 331454 262734 331538
rect 262114 331218 262146 331454
rect 262382 331218 262466 331454
rect 262702 331218 262734 331454
rect 262114 297774 262734 331218
rect 262114 297538 262146 297774
rect 262382 297538 262466 297774
rect 262702 297538 262734 297774
rect 262114 297454 262734 297538
rect 262114 297218 262146 297454
rect 262382 297218 262466 297454
rect 262702 297218 262734 297454
rect 262114 263774 262734 297218
rect 262114 263538 262146 263774
rect 262382 263538 262466 263774
rect 262702 263538 262734 263774
rect 262114 263454 262734 263538
rect 262114 263218 262146 263454
rect 262382 263218 262466 263454
rect 262702 263218 262734 263454
rect 262114 229774 262734 263218
rect 262114 229538 262146 229774
rect 262382 229538 262466 229774
rect 262702 229538 262734 229774
rect 262114 229454 262734 229538
rect 262114 229218 262146 229454
rect 262382 229218 262466 229454
rect 262702 229218 262734 229454
rect 262114 225660 262734 229218
rect 265834 711558 266454 711590
rect 265834 711322 265866 711558
rect 266102 711322 266186 711558
rect 266422 711322 266454 711558
rect 265834 711238 266454 711322
rect 265834 711002 265866 711238
rect 266102 711002 266186 711238
rect 266422 711002 266454 711238
rect 265834 675494 266454 711002
rect 265834 675258 265866 675494
rect 266102 675258 266186 675494
rect 266422 675258 266454 675494
rect 265834 675174 266454 675258
rect 265834 674938 265866 675174
rect 266102 674938 266186 675174
rect 266422 674938 266454 675174
rect 265834 641494 266454 674938
rect 265834 641258 265866 641494
rect 266102 641258 266186 641494
rect 266422 641258 266454 641494
rect 265834 641174 266454 641258
rect 265834 640938 265866 641174
rect 266102 640938 266186 641174
rect 266422 640938 266454 641174
rect 265834 607494 266454 640938
rect 265834 607258 265866 607494
rect 266102 607258 266186 607494
rect 266422 607258 266454 607494
rect 265834 607174 266454 607258
rect 265834 606938 265866 607174
rect 266102 606938 266186 607174
rect 266422 606938 266454 607174
rect 265834 573494 266454 606938
rect 265834 573258 265866 573494
rect 266102 573258 266186 573494
rect 266422 573258 266454 573494
rect 265834 573174 266454 573258
rect 265834 572938 265866 573174
rect 266102 572938 266186 573174
rect 266422 572938 266454 573174
rect 265834 539494 266454 572938
rect 265834 539258 265866 539494
rect 266102 539258 266186 539494
rect 266422 539258 266454 539494
rect 265834 539174 266454 539258
rect 265834 538938 265866 539174
rect 266102 538938 266186 539174
rect 266422 538938 266454 539174
rect 265834 505494 266454 538938
rect 265834 505258 265866 505494
rect 266102 505258 266186 505494
rect 266422 505258 266454 505494
rect 265834 505174 266454 505258
rect 265834 504938 265866 505174
rect 266102 504938 266186 505174
rect 266422 504938 266454 505174
rect 265834 471494 266454 504938
rect 265834 471258 265866 471494
rect 266102 471258 266186 471494
rect 266422 471258 266454 471494
rect 265834 471174 266454 471258
rect 265834 470938 265866 471174
rect 266102 470938 266186 471174
rect 266422 470938 266454 471174
rect 265834 437494 266454 470938
rect 265834 437258 265866 437494
rect 266102 437258 266186 437494
rect 266422 437258 266454 437494
rect 265834 437174 266454 437258
rect 265834 436938 265866 437174
rect 266102 436938 266186 437174
rect 266422 436938 266454 437174
rect 265834 403494 266454 436938
rect 265834 403258 265866 403494
rect 266102 403258 266186 403494
rect 266422 403258 266454 403494
rect 265834 403174 266454 403258
rect 265834 402938 265866 403174
rect 266102 402938 266186 403174
rect 266422 402938 266454 403174
rect 265834 369494 266454 402938
rect 265834 369258 265866 369494
rect 266102 369258 266186 369494
rect 266422 369258 266454 369494
rect 265834 369174 266454 369258
rect 265834 368938 265866 369174
rect 266102 368938 266186 369174
rect 266422 368938 266454 369174
rect 265834 335494 266454 368938
rect 265834 335258 265866 335494
rect 266102 335258 266186 335494
rect 266422 335258 266454 335494
rect 265834 335174 266454 335258
rect 265834 334938 265866 335174
rect 266102 334938 266186 335174
rect 266422 334938 266454 335174
rect 265834 301494 266454 334938
rect 265834 301258 265866 301494
rect 266102 301258 266186 301494
rect 266422 301258 266454 301494
rect 265834 301174 266454 301258
rect 265834 300938 265866 301174
rect 266102 300938 266186 301174
rect 266422 300938 266454 301174
rect 265834 267494 266454 300938
rect 265834 267258 265866 267494
rect 266102 267258 266186 267494
rect 266422 267258 266454 267494
rect 265834 267174 266454 267258
rect 265834 266938 265866 267174
rect 266102 266938 266186 267174
rect 266422 266938 266454 267174
rect 265834 233494 266454 266938
rect 265834 233258 265866 233494
rect 266102 233258 266186 233494
rect 266422 233258 266454 233494
rect 265834 233174 266454 233258
rect 265834 232938 265866 233174
rect 266102 232938 266186 233174
rect 266422 232938 266454 233174
rect 265834 225660 266454 232938
rect 273794 704838 274414 711590
rect 273794 704602 273826 704838
rect 274062 704602 274146 704838
rect 274382 704602 274414 704838
rect 273794 704518 274414 704602
rect 273794 704282 273826 704518
rect 274062 704282 274146 704518
rect 274382 704282 274414 704518
rect 273794 683454 274414 704282
rect 273794 683218 273826 683454
rect 274062 683218 274146 683454
rect 274382 683218 274414 683454
rect 273794 683134 274414 683218
rect 273794 682898 273826 683134
rect 274062 682898 274146 683134
rect 274382 682898 274414 683134
rect 273794 649454 274414 682898
rect 273794 649218 273826 649454
rect 274062 649218 274146 649454
rect 274382 649218 274414 649454
rect 273794 649134 274414 649218
rect 273794 648898 273826 649134
rect 274062 648898 274146 649134
rect 274382 648898 274414 649134
rect 273794 615454 274414 648898
rect 273794 615218 273826 615454
rect 274062 615218 274146 615454
rect 274382 615218 274414 615454
rect 273794 615134 274414 615218
rect 273794 614898 273826 615134
rect 274062 614898 274146 615134
rect 274382 614898 274414 615134
rect 273794 581454 274414 614898
rect 273794 581218 273826 581454
rect 274062 581218 274146 581454
rect 274382 581218 274414 581454
rect 273794 581134 274414 581218
rect 273794 580898 273826 581134
rect 274062 580898 274146 581134
rect 274382 580898 274414 581134
rect 273794 547454 274414 580898
rect 273794 547218 273826 547454
rect 274062 547218 274146 547454
rect 274382 547218 274414 547454
rect 273794 547134 274414 547218
rect 273794 546898 273826 547134
rect 274062 546898 274146 547134
rect 274382 546898 274414 547134
rect 273794 513454 274414 546898
rect 273794 513218 273826 513454
rect 274062 513218 274146 513454
rect 274382 513218 274414 513454
rect 273794 513134 274414 513218
rect 273794 512898 273826 513134
rect 274062 512898 274146 513134
rect 274382 512898 274414 513134
rect 273794 479454 274414 512898
rect 273794 479218 273826 479454
rect 274062 479218 274146 479454
rect 274382 479218 274414 479454
rect 273794 479134 274414 479218
rect 273794 478898 273826 479134
rect 274062 478898 274146 479134
rect 274382 478898 274414 479134
rect 273794 445454 274414 478898
rect 273794 445218 273826 445454
rect 274062 445218 274146 445454
rect 274382 445218 274414 445454
rect 273794 445134 274414 445218
rect 273794 444898 273826 445134
rect 274062 444898 274146 445134
rect 274382 444898 274414 445134
rect 273794 411454 274414 444898
rect 273794 411218 273826 411454
rect 274062 411218 274146 411454
rect 274382 411218 274414 411454
rect 273794 411134 274414 411218
rect 273794 410898 273826 411134
rect 274062 410898 274146 411134
rect 274382 410898 274414 411134
rect 273794 377454 274414 410898
rect 273794 377218 273826 377454
rect 274062 377218 274146 377454
rect 274382 377218 274414 377454
rect 273794 377134 274414 377218
rect 273794 376898 273826 377134
rect 274062 376898 274146 377134
rect 274382 376898 274414 377134
rect 273794 343454 274414 376898
rect 273794 343218 273826 343454
rect 274062 343218 274146 343454
rect 274382 343218 274414 343454
rect 273794 343134 274414 343218
rect 273794 342898 273826 343134
rect 274062 342898 274146 343134
rect 274382 342898 274414 343134
rect 273794 309454 274414 342898
rect 273794 309218 273826 309454
rect 274062 309218 274146 309454
rect 274382 309218 274414 309454
rect 273794 309134 274414 309218
rect 273794 308898 273826 309134
rect 274062 308898 274146 309134
rect 274382 308898 274414 309134
rect 273794 275454 274414 308898
rect 273794 275218 273826 275454
rect 274062 275218 274146 275454
rect 274382 275218 274414 275454
rect 273794 275134 274414 275218
rect 273794 274898 273826 275134
rect 274062 274898 274146 275134
rect 274382 274898 274414 275134
rect 273794 241454 274414 274898
rect 273794 241218 273826 241454
rect 274062 241218 274146 241454
rect 274382 241218 274414 241454
rect 273794 241134 274414 241218
rect 273794 240898 273826 241134
rect 274062 240898 274146 241134
rect 274382 240898 274414 241134
rect 273794 225660 274414 240898
rect 277514 705798 278134 711590
rect 277514 705562 277546 705798
rect 277782 705562 277866 705798
rect 278102 705562 278134 705798
rect 277514 705478 278134 705562
rect 277514 705242 277546 705478
rect 277782 705242 277866 705478
rect 278102 705242 278134 705478
rect 277514 687174 278134 705242
rect 277514 686938 277546 687174
rect 277782 686938 277866 687174
rect 278102 686938 278134 687174
rect 277514 686854 278134 686938
rect 277514 686618 277546 686854
rect 277782 686618 277866 686854
rect 278102 686618 278134 686854
rect 277514 653174 278134 686618
rect 277514 652938 277546 653174
rect 277782 652938 277866 653174
rect 278102 652938 278134 653174
rect 277514 652854 278134 652938
rect 277514 652618 277546 652854
rect 277782 652618 277866 652854
rect 278102 652618 278134 652854
rect 277514 619174 278134 652618
rect 277514 618938 277546 619174
rect 277782 618938 277866 619174
rect 278102 618938 278134 619174
rect 277514 618854 278134 618938
rect 277514 618618 277546 618854
rect 277782 618618 277866 618854
rect 278102 618618 278134 618854
rect 277514 585174 278134 618618
rect 277514 584938 277546 585174
rect 277782 584938 277866 585174
rect 278102 584938 278134 585174
rect 277514 584854 278134 584938
rect 277514 584618 277546 584854
rect 277782 584618 277866 584854
rect 278102 584618 278134 584854
rect 277514 551174 278134 584618
rect 277514 550938 277546 551174
rect 277782 550938 277866 551174
rect 278102 550938 278134 551174
rect 277514 550854 278134 550938
rect 277514 550618 277546 550854
rect 277782 550618 277866 550854
rect 278102 550618 278134 550854
rect 277514 517174 278134 550618
rect 277514 516938 277546 517174
rect 277782 516938 277866 517174
rect 278102 516938 278134 517174
rect 277514 516854 278134 516938
rect 277514 516618 277546 516854
rect 277782 516618 277866 516854
rect 278102 516618 278134 516854
rect 277514 483174 278134 516618
rect 277514 482938 277546 483174
rect 277782 482938 277866 483174
rect 278102 482938 278134 483174
rect 277514 482854 278134 482938
rect 277514 482618 277546 482854
rect 277782 482618 277866 482854
rect 278102 482618 278134 482854
rect 277514 449174 278134 482618
rect 277514 448938 277546 449174
rect 277782 448938 277866 449174
rect 278102 448938 278134 449174
rect 277514 448854 278134 448938
rect 277514 448618 277546 448854
rect 277782 448618 277866 448854
rect 278102 448618 278134 448854
rect 277514 415174 278134 448618
rect 277514 414938 277546 415174
rect 277782 414938 277866 415174
rect 278102 414938 278134 415174
rect 277514 414854 278134 414938
rect 277514 414618 277546 414854
rect 277782 414618 277866 414854
rect 278102 414618 278134 414854
rect 277514 381174 278134 414618
rect 277514 380938 277546 381174
rect 277782 380938 277866 381174
rect 278102 380938 278134 381174
rect 277514 380854 278134 380938
rect 277514 380618 277546 380854
rect 277782 380618 277866 380854
rect 278102 380618 278134 380854
rect 277514 347174 278134 380618
rect 277514 346938 277546 347174
rect 277782 346938 277866 347174
rect 278102 346938 278134 347174
rect 277514 346854 278134 346938
rect 277514 346618 277546 346854
rect 277782 346618 277866 346854
rect 278102 346618 278134 346854
rect 277514 313174 278134 346618
rect 277514 312938 277546 313174
rect 277782 312938 277866 313174
rect 278102 312938 278134 313174
rect 277514 312854 278134 312938
rect 277514 312618 277546 312854
rect 277782 312618 277866 312854
rect 278102 312618 278134 312854
rect 277514 279174 278134 312618
rect 277514 278938 277546 279174
rect 277782 278938 277866 279174
rect 278102 278938 278134 279174
rect 277514 278854 278134 278938
rect 277514 278618 277546 278854
rect 277782 278618 277866 278854
rect 278102 278618 278134 278854
rect 277514 245174 278134 278618
rect 277514 244938 277546 245174
rect 277782 244938 277866 245174
rect 278102 244938 278134 245174
rect 277514 244854 278134 244938
rect 277514 244618 277546 244854
rect 277782 244618 277866 244854
rect 278102 244618 278134 244854
rect 277514 225660 278134 244618
rect 281234 706758 281854 711590
rect 281234 706522 281266 706758
rect 281502 706522 281586 706758
rect 281822 706522 281854 706758
rect 281234 706438 281854 706522
rect 281234 706202 281266 706438
rect 281502 706202 281586 706438
rect 281822 706202 281854 706438
rect 281234 690894 281854 706202
rect 281234 690658 281266 690894
rect 281502 690658 281586 690894
rect 281822 690658 281854 690894
rect 281234 690574 281854 690658
rect 281234 690338 281266 690574
rect 281502 690338 281586 690574
rect 281822 690338 281854 690574
rect 281234 656894 281854 690338
rect 281234 656658 281266 656894
rect 281502 656658 281586 656894
rect 281822 656658 281854 656894
rect 281234 656574 281854 656658
rect 281234 656338 281266 656574
rect 281502 656338 281586 656574
rect 281822 656338 281854 656574
rect 281234 622894 281854 656338
rect 281234 622658 281266 622894
rect 281502 622658 281586 622894
rect 281822 622658 281854 622894
rect 281234 622574 281854 622658
rect 281234 622338 281266 622574
rect 281502 622338 281586 622574
rect 281822 622338 281854 622574
rect 281234 588894 281854 622338
rect 281234 588658 281266 588894
rect 281502 588658 281586 588894
rect 281822 588658 281854 588894
rect 281234 588574 281854 588658
rect 281234 588338 281266 588574
rect 281502 588338 281586 588574
rect 281822 588338 281854 588574
rect 281234 554894 281854 588338
rect 281234 554658 281266 554894
rect 281502 554658 281586 554894
rect 281822 554658 281854 554894
rect 281234 554574 281854 554658
rect 281234 554338 281266 554574
rect 281502 554338 281586 554574
rect 281822 554338 281854 554574
rect 281234 520894 281854 554338
rect 281234 520658 281266 520894
rect 281502 520658 281586 520894
rect 281822 520658 281854 520894
rect 281234 520574 281854 520658
rect 281234 520338 281266 520574
rect 281502 520338 281586 520574
rect 281822 520338 281854 520574
rect 281234 486894 281854 520338
rect 281234 486658 281266 486894
rect 281502 486658 281586 486894
rect 281822 486658 281854 486894
rect 281234 486574 281854 486658
rect 281234 486338 281266 486574
rect 281502 486338 281586 486574
rect 281822 486338 281854 486574
rect 281234 452894 281854 486338
rect 281234 452658 281266 452894
rect 281502 452658 281586 452894
rect 281822 452658 281854 452894
rect 281234 452574 281854 452658
rect 281234 452338 281266 452574
rect 281502 452338 281586 452574
rect 281822 452338 281854 452574
rect 281234 418894 281854 452338
rect 281234 418658 281266 418894
rect 281502 418658 281586 418894
rect 281822 418658 281854 418894
rect 281234 418574 281854 418658
rect 281234 418338 281266 418574
rect 281502 418338 281586 418574
rect 281822 418338 281854 418574
rect 281234 384894 281854 418338
rect 281234 384658 281266 384894
rect 281502 384658 281586 384894
rect 281822 384658 281854 384894
rect 281234 384574 281854 384658
rect 281234 384338 281266 384574
rect 281502 384338 281586 384574
rect 281822 384338 281854 384574
rect 281234 350894 281854 384338
rect 281234 350658 281266 350894
rect 281502 350658 281586 350894
rect 281822 350658 281854 350894
rect 281234 350574 281854 350658
rect 281234 350338 281266 350574
rect 281502 350338 281586 350574
rect 281822 350338 281854 350574
rect 281234 316894 281854 350338
rect 281234 316658 281266 316894
rect 281502 316658 281586 316894
rect 281822 316658 281854 316894
rect 281234 316574 281854 316658
rect 281234 316338 281266 316574
rect 281502 316338 281586 316574
rect 281822 316338 281854 316574
rect 281234 282894 281854 316338
rect 281234 282658 281266 282894
rect 281502 282658 281586 282894
rect 281822 282658 281854 282894
rect 281234 282574 281854 282658
rect 281234 282338 281266 282574
rect 281502 282338 281586 282574
rect 281822 282338 281854 282574
rect 281234 248894 281854 282338
rect 281234 248658 281266 248894
rect 281502 248658 281586 248894
rect 281822 248658 281854 248894
rect 281234 248574 281854 248658
rect 281234 248338 281266 248574
rect 281502 248338 281586 248574
rect 281822 248338 281854 248574
rect 250954 218378 250986 218614
rect 251222 218378 251306 218614
rect 251542 218378 251574 218614
rect 250954 218294 251574 218378
rect 250954 218058 250986 218294
rect 251222 218058 251306 218294
rect 251542 218058 251574 218294
rect 220674 188098 220706 188334
rect 220942 188098 221026 188334
rect 221262 188098 221294 188334
rect 220674 188014 221294 188098
rect 220674 187778 220706 188014
rect 220942 187778 221026 188014
rect 221262 187778 221294 188014
rect 220674 154334 221294 187778
rect 220674 154098 220706 154334
rect 220942 154098 221026 154334
rect 221262 154098 221294 154334
rect 220674 154014 221294 154098
rect 220674 153778 220706 154014
rect 220942 153778 221026 154014
rect 221262 153778 221294 154014
rect 220674 120334 221294 153778
rect 220674 120098 220706 120334
rect 220942 120098 221026 120334
rect 221262 120098 221294 120334
rect 220674 120014 221294 120098
rect 220674 119778 220706 120014
rect 220942 119778 221026 120014
rect 221262 119778 221294 120014
rect 220674 86334 221294 119778
rect 220674 86098 220706 86334
rect 220942 86098 221026 86334
rect 221262 86098 221294 86334
rect 220674 86014 221294 86098
rect 220674 85778 220706 86014
rect 220942 85778 221026 86014
rect 221262 85778 221294 86014
rect 220674 52334 221294 85778
rect 220674 52098 220706 52334
rect 220942 52098 221026 52334
rect 221262 52098 221294 52334
rect 220674 52014 221294 52098
rect 220674 51778 220706 52014
rect 220942 51778 221026 52014
rect 221262 51778 221294 52014
rect 220674 18334 221294 51778
rect 220674 18098 220706 18334
rect 220942 18098 221026 18334
rect 221262 18098 221294 18334
rect 220674 18014 221294 18098
rect 220674 17778 220706 18014
rect 220942 17778 221026 18014
rect 221262 17778 221294 18014
rect 220674 -4186 221294 17778
rect 220674 -4422 220706 -4186
rect 220942 -4422 221026 -4186
rect 221262 -4422 221294 -4186
rect 220674 -4506 221294 -4422
rect 220674 -4742 220706 -4506
rect 220942 -4742 221026 -4506
rect 221262 -4742 221294 -4506
rect 220674 -7654 221294 -4742
rect 224394 192054 225014 214340
rect 224394 191818 224426 192054
rect 224662 191818 224746 192054
rect 224982 191818 225014 192054
rect 224394 191734 225014 191818
rect 224394 191498 224426 191734
rect 224662 191498 224746 191734
rect 224982 191498 225014 191734
rect 224394 158054 225014 191498
rect 224394 157818 224426 158054
rect 224662 157818 224746 158054
rect 224982 157818 225014 158054
rect 224394 157734 225014 157818
rect 224394 157498 224426 157734
rect 224662 157498 224746 157734
rect 224982 157498 225014 157734
rect 224394 124054 225014 157498
rect 224394 123818 224426 124054
rect 224662 123818 224746 124054
rect 224982 123818 225014 124054
rect 224394 123734 225014 123818
rect 224394 123498 224426 123734
rect 224662 123498 224746 123734
rect 224982 123498 225014 123734
rect 224394 90054 225014 123498
rect 224394 89818 224426 90054
rect 224662 89818 224746 90054
rect 224982 89818 225014 90054
rect 224394 89734 225014 89818
rect 224394 89498 224426 89734
rect 224662 89498 224746 89734
rect 224982 89498 225014 89734
rect 224394 56054 225014 89498
rect 224394 55818 224426 56054
rect 224662 55818 224746 56054
rect 224982 55818 225014 56054
rect 224394 55734 225014 55818
rect 224394 55498 224426 55734
rect 224662 55498 224746 55734
rect 224982 55498 225014 55734
rect 224394 22054 225014 55498
rect 224394 21818 224426 22054
rect 224662 21818 224746 22054
rect 224982 21818 225014 22054
rect 224394 21734 225014 21818
rect 224394 21498 224426 21734
rect 224662 21498 224746 21734
rect 224982 21498 225014 21734
rect 224394 -5146 225014 21498
rect 224394 -5382 224426 -5146
rect 224662 -5382 224746 -5146
rect 224982 -5382 225014 -5146
rect 224394 -5466 225014 -5382
rect 224394 -5702 224426 -5466
rect 224662 -5702 224746 -5466
rect 224982 -5702 225014 -5466
rect 224394 -7654 225014 -5702
rect 228114 195774 228734 214340
rect 228114 195538 228146 195774
rect 228382 195538 228466 195774
rect 228702 195538 228734 195774
rect 228114 195454 228734 195538
rect 228114 195218 228146 195454
rect 228382 195218 228466 195454
rect 228702 195218 228734 195454
rect 228114 161774 228734 195218
rect 228114 161538 228146 161774
rect 228382 161538 228466 161774
rect 228702 161538 228734 161774
rect 228114 161454 228734 161538
rect 228114 161218 228146 161454
rect 228382 161218 228466 161454
rect 228702 161218 228734 161454
rect 228114 127774 228734 161218
rect 228114 127538 228146 127774
rect 228382 127538 228466 127774
rect 228702 127538 228734 127774
rect 228114 127454 228734 127538
rect 228114 127218 228146 127454
rect 228382 127218 228466 127454
rect 228702 127218 228734 127454
rect 228114 93774 228734 127218
rect 228114 93538 228146 93774
rect 228382 93538 228466 93774
rect 228702 93538 228734 93774
rect 228114 93454 228734 93538
rect 228114 93218 228146 93454
rect 228382 93218 228466 93454
rect 228702 93218 228734 93454
rect 228114 59774 228734 93218
rect 228114 59538 228146 59774
rect 228382 59538 228466 59774
rect 228702 59538 228734 59774
rect 228114 59454 228734 59538
rect 228114 59218 228146 59454
rect 228382 59218 228466 59454
rect 228702 59218 228734 59454
rect 228114 25774 228734 59218
rect 228114 25538 228146 25774
rect 228382 25538 228466 25774
rect 228702 25538 228734 25774
rect 228114 25454 228734 25538
rect 228114 25218 228146 25454
rect 228382 25218 228466 25454
rect 228702 25218 228734 25454
rect 228114 -6106 228734 25218
rect 228114 -6342 228146 -6106
rect 228382 -6342 228466 -6106
rect 228702 -6342 228734 -6106
rect 228114 -6426 228734 -6342
rect 228114 -6662 228146 -6426
rect 228382 -6662 228466 -6426
rect 228702 -6662 228734 -6426
rect 228114 -7654 228734 -6662
rect 231834 199494 232454 214340
rect 231834 199258 231866 199494
rect 232102 199258 232186 199494
rect 232422 199258 232454 199494
rect 231834 199174 232454 199258
rect 231834 198938 231866 199174
rect 232102 198938 232186 199174
rect 232422 198938 232454 199174
rect 231834 165494 232454 198938
rect 231834 165258 231866 165494
rect 232102 165258 232186 165494
rect 232422 165258 232454 165494
rect 231834 165174 232454 165258
rect 231834 164938 231866 165174
rect 232102 164938 232186 165174
rect 232422 164938 232454 165174
rect 231834 131494 232454 164938
rect 231834 131258 231866 131494
rect 232102 131258 232186 131494
rect 232422 131258 232454 131494
rect 231834 131174 232454 131258
rect 231834 130938 231866 131174
rect 232102 130938 232186 131174
rect 232422 130938 232454 131174
rect 231834 97494 232454 130938
rect 231834 97258 231866 97494
rect 232102 97258 232186 97494
rect 232422 97258 232454 97494
rect 231834 97174 232454 97258
rect 231834 96938 231866 97174
rect 232102 96938 232186 97174
rect 232422 96938 232454 97174
rect 231834 63494 232454 96938
rect 231834 63258 231866 63494
rect 232102 63258 232186 63494
rect 232422 63258 232454 63494
rect 231834 63174 232454 63258
rect 231834 62938 231866 63174
rect 232102 62938 232186 63174
rect 232422 62938 232454 63174
rect 231834 29494 232454 62938
rect 231834 29258 231866 29494
rect 232102 29258 232186 29494
rect 232422 29258 232454 29494
rect 231834 29174 232454 29258
rect 231834 28938 231866 29174
rect 232102 28938 232186 29174
rect 232422 28938 232454 29174
rect 231834 -7066 232454 28938
rect 231834 -7302 231866 -7066
rect 232102 -7302 232186 -7066
rect 232422 -7302 232454 -7066
rect 231834 -7386 232454 -7302
rect 231834 -7622 231866 -7386
rect 232102 -7622 232186 -7386
rect 232422 -7622 232454 -7386
rect 231834 -7654 232454 -7622
rect 239794 207454 240414 214340
rect 239794 207218 239826 207454
rect 240062 207218 240146 207454
rect 240382 207218 240414 207454
rect 239794 207134 240414 207218
rect 239794 206898 239826 207134
rect 240062 206898 240146 207134
rect 240382 206898 240414 207134
rect 239794 173454 240414 206898
rect 239794 173218 239826 173454
rect 240062 173218 240146 173454
rect 240382 173218 240414 173454
rect 239794 173134 240414 173218
rect 239794 172898 239826 173134
rect 240062 172898 240146 173134
rect 240382 172898 240414 173134
rect 239794 139454 240414 172898
rect 239794 139218 239826 139454
rect 240062 139218 240146 139454
rect 240382 139218 240414 139454
rect 239794 139134 240414 139218
rect 239794 138898 239826 139134
rect 240062 138898 240146 139134
rect 240382 138898 240414 139134
rect 239794 105454 240414 138898
rect 239794 105218 239826 105454
rect 240062 105218 240146 105454
rect 240382 105218 240414 105454
rect 239794 105134 240414 105218
rect 239794 104898 239826 105134
rect 240062 104898 240146 105134
rect 240382 104898 240414 105134
rect 239794 71454 240414 104898
rect 239794 71218 239826 71454
rect 240062 71218 240146 71454
rect 240382 71218 240414 71454
rect 239794 71134 240414 71218
rect 239794 70898 239826 71134
rect 240062 70898 240146 71134
rect 240382 70898 240414 71134
rect 239794 37454 240414 70898
rect 239794 37218 239826 37454
rect 240062 37218 240146 37454
rect 240382 37218 240414 37454
rect 239794 37134 240414 37218
rect 239794 36898 239826 37134
rect 240062 36898 240146 37134
rect 240382 36898 240414 37134
rect 239794 3454 240414 36898
rect 239794 3218 239826 3454
rect 240062 3218 240146 3454
rect 240382 3218 240414 3454
rect 239794 3134 240414 3218
rect 239794 2898 239826 3134
rect 240062 2898 240146 3134
rect 240382 2898 240414 3134
rect 239794 -346 240414 2898
rect 239794 -582 239826 -346
rect 240062 -582 240146 -346
rect 240382 -582 240414 -346
rect 239794 -666 240414 -582
rect 239794 -902 239826 -666
rect 240062 -902 240146 -666
rect 240382 -902 240414 -666
rect 239794 -7654 240414 -902
rect 243514 211174 244134 214340
rect 243514 210938 243546 211174
rect 243782 210938 243866 211174
rect 244102 210938 244134 211174
rect 243514 210854 244134 210938
rect 243514 210618 243546 210854
rect 243782 210618 243866 210854
rect 244102 210618 244134 210854
rect 243514 177174 244134 210618
rect 243514 176938 243546 177174
rect 243782 176938 243866 177174
rect 244102 176938 244134 177174
rect 243514 176854 244134 176938
rect 243514 176618 243546 176854
rect 243782 176618 243866 176854
rect 244102 176618 244134 176854
rect 243514 143174 244134 176618
rect 243514 142938 243546 143174
rect 243782 142938 243866 143174
rect 244102 142938 244134 143174
rect 243514 142854 244134 142938
rect 243514 142618 243546 142854
rect 243782 142618 243866 142854
rect 244102 142618 244134 142854
rect 243514 109174 244134 142618
rect 243514 108938 243546 109174
rect 243782 108938 243866 109174
rect 244102 108938 244134 109174
rect 243514 108854 244134 108938
rect 243514 108618 243546 108854
rect 243782 108618 243866 108854
rect 244102 108618 244134 108854
rect 243514 75174 244134 108618
rect 243514 74938 243546 75174
rect 243782 74938 243866 75174
rect 244102 74938 244134 75174
rect 243514 74854 244134 74938
rect 243514 74618 243546 74854
rect 243782 74618 243866 74854
rect 244102 74618 244134 74854
rect 243514 41174 244134 74618
rect 243514 40938 243546 41174
rect 243782 40938 243866 41174
rect 244102 40938 244134 41174
rect 243514 40854 244134 40938
rect 243514 40618 243546 40854
rect 243782 40618 243866 40854
rect 244102 40618 244134 40854
rect 243514 7174 244134 40618
rect 243514 6938 243546 7174
rect 243782 6938 243866 7174
rect 244102 6938 244134 7174
rect 243514 6854 244134 6938
rect 243514 6618 243546 6854
rect 243782 6618 243866 6854
rect 244102 6618 244134 6854
rect 243514 -1306 244134 6618
rect 243514 -1542 243546 -1306
rect 243782 -1542 243866 -1306
rect 244102 -1542 244134 -1306
rect 243514 -1626 244134 -1542
rect 243514 -1862 243546 -1626
rect 243782 -1862 243866 -1626
rect 244102 -1862 244134 -1626
rect 243514 -7654 244134 -1862
rect 247234 180894 247854 214340
rect 247234 180658 247266 180894
rect 247502 180658 247586 180894
rect 247822 180658 247854 180894
rect 247234 180574 247854 180658
rect 247234 180338 247266 180574
rect 247502 180338 247586 180574
rect 247822 180338 247854 180574
rect 247234 146894 247854 180338
rect 247234 146658 247266 146894
rect 247502 146658 247586 146894
rect 247822 146658 247854 146894
rect 247234 146574 247854 146658
rect 247234 146338 247266 146574
rect 247502 146338 247586 146574
rect 247822 146338 247854 146574
rect 247234 112894 247854 146338
rect 247234 112658 247266 112894
rect 247502 112658 247586 112894
rect 247822 112658 247854 112894
rect 247234 112574 247854 112658
rect 247234 112338 247266 112574
rect 247502 112338 247586 112574
rect 247822 112338 247854 112574
rect 247234 78894 247854 112338
rect 247234 78658 247266 78894
rect 247502 78658 247586 78894
rect 247822 78658 247854 78894
rect 247234 78574 247854 78658
rect 247234 78338 247266 78574
rect 247502 78338 247586 78574
rect 247822 78338 247854 78574
rect 247234 44894 247854 78338
rect 247234 44658 247266 44894
rect 247502 44658 247586 44894
rect 247822 44658 247854 44894
rect 247234 44574 247854 44658
rect 247234 44338 247266 44574
rect 247502 44338 247586 44574
rect 247822 44338 247854 44574
rect 247234 10894 247854 44338
rect 247234 10658 247266 10894
rect 247502 10658 247586 10894
rect 247822 10658 247854 10894
rect 247234 10574 247854 10658
rect 247234 10338 247266 10574
rect 247502 10338 247586 10574
rect 247822 10338 247854 10574
rect 247234 -2266 247854 10338
rect 247234 -2502 247266 -2266
rect 247502 -2502 247586 -2266
rect 247822 -2502 247854 -2266
rect 247234 -2586 247854 -2502
rect 247234 -2822 247266 -2586
rect 247502 -2822 247586 -2586
rect 247822 -2822 247854 -2586
rect 247234 -7654 247854 -2822
rect 250954 184614 251574 218058
rect 281234 214894 281854 248338
rect 284954 707718 285574 711590
rect 284954 707482 284986 707718
rect 285222 707482 285306 707718
rect 285542 707482 285574 707718
rect 284954 707398 285574 707482
rect 284954 707162 284986 707398
rect 285222 707162 285306 707398
rect 285542 707162 285574 707398
rect 284954 694614 285574 707162
rect 284954 694378 284986 694614
rect 285222 694378 285306 694614
rect 285542 694378 285574 694614
rect 284954 694294 285574 694378
rect 284954 694058 284986 694294
rect 285222 694058 285306 694294
rect 285542 694058 285574 694294
rect 284954 660614 285574 694058
rect 284954 660378 284986 660614
rect 285222 660378 285306 660614
rect 285542 660378 285574 660614
rect 284954 660294 285574 660378
rect 284954 660058 284986 660294
rect 285222 660058 285306 660294
rect 285542 660058 285574 660294
rect 284954 626614 285574 660058
rect 284954 626378 284986 626614
rect 285222 626378 285306 626614
rect 285542 626378 285574 626614
rect 284954 626294 285574 626378
rect 284954 626058 284986 626294
rect 285222 626058 285306 626294
rect 285542 626058 285574 626294
rect 284954 592614 285574 626058
rect 284954 592378 284986 592614
rect 285222 592378 285306 592614
rect 285542 592378 285574 592614
rect 284954 592294 285574 592378
rect 284954 592058 284986 592294
rect 285222 592058 285306 592294
rect 285542 592058 285574 592294
rect 284954 558614 285574 592058
rect 284954 558378 284986 558614
rect 285222 558378 285306 558614
rect 285542 558378 285574 558614
rect 284954 558294 285574 558378
rect 284954 558058 284986 558294
rect 285222 558058 285306 558294
rect 285542 558058 285574 558294
rect 284954 524614 285574 558058
rect 284954 524378 284986 524614
rect 285222 524378 285306 524614
rect 285542 524378 285574 524614
rect 284954 524294 285574 524378
rect 284954 524058 284986 524294
rect 285222 524058 285306 524294
rect 285542 524058 285574 524294
rect 284954 490614 285574 524058
rect 284954 490378 284986 490614
rect 285222 490378 285306 490614
rect 285542 490378 285574 490614
rect 284954 490294 285574 490378
rect 284954 490058 284986 490294
rect 285222 490058 285306 490294
rect 285542 490058 285574 490294
rect 284954 456614 285574 490058
rect 284954 456378 284986 456614
rect 285222 456378 285306 456614
rect 285542 456378 285574 456614
rect 284954 456294 285574 456378
rect 284954 456058 284986 456294
rect 285222 456058 285306 456294
rect 285542 456058 285574 456294
rect 284954 422614 285574 456058
rect 284954 422378 284986 422614
rect 285222 422378 285306 422614
rect 285542 422378 285574 422614
rect 284954 422294 285574 422378
rect 284954 422058 284986 422294
rect 285222 422058 285306 422294
rect 285542 422058 285574 422294
rect 284954 388614 285574 422058
rect 284954 388378 284986 388614
rect 285222 388378 285306 388614
rect 285542 388378 285574 388614
rect 284954 388294 285574 388378
rect 284954 388058 284986 388294
rect 285222 388058 285306 388294
rect 285542 388058 285574 388294
rect 284954 354614 285574 388058
rect 284954 354378 284986 354614
rect 285222 354378 285306 354614
rect 285542 354378 285574 354614
rect 284954 354294 285574 354378
rect 284954 354058 284986 354294
rect 285222 354058 285306 354294
rect 285542 354058 285574 354294
rect 284954 320614 285574 354058
rect 284954 320378 284986 320614
rect 285222 320378 285306 320614
rect 285542 320378 285574 320614
rect 284954 320294 285574 320378
rect 284954 320058 284986 320294
rect 285222 320058 285306 320294
rect 285542 320058 285574 320294
rect 284954 286614 285574 320058
rect 284954 286378 284986 286614
rect 285222 286378 285306 286614
rect 285542 286378 285574 286614
rect 284954 286294 285574 286378
rect 284954 286058 284986 286294
rect 285222 286058 285306 286294
rect 285542 286058 285574 286294
rect 284954 252614 285574 286058
rect 284954 252378 284986 252614
rect 285222 252378 285306 252614
rect 285542 252378 285574 252614
rect 284954 252294 285574 252378
rect 284954 252058 284986 252294
rect 285222 252058 285306 252294
rect 285542 252058 285574 252294
rect 284954 225660 285574 252058
rect 288674 708678 289294 711590
rect 288674 708442 288706 708678
rect 288942 708442 289026 708678
rect 289262 708442 289294 708678
rect 288674 708358 289294 708442
rect 288674 708122 288706 708358
rect 288942 708122 289026 708358
rect 289262 708122 289294 708358
rect 288674 698334 289294 708122
rect 288674 698098 288706 698334
rect 288942 698098 289026 698334
rect 289262 698098 289294 698334
rect 288674 698014 289294 698098
rect 288674 697778 288706 698014
rect 288942 697778 289026 698014
rect 289262 697778 289294 698014
rect 288674 664334 289294 697778
rect 288674 664098 288706 664334
rect 288942 664098 289026 664334
rect 289262 664098 289294 664334
rect 288674 664014 289294 664098
rect 288674 663778 288706 664014
rect 288942 663778 289026 664014
rect 289262 663778 289294 664014
rect 288674 630334 289294 663778
rect 288674 630098 288706 630334
rect 288942 630098 289026 630334
rect 289262 630098 289294 630334
rect 288674 630014 289294 630098
rect 288674 629778 288706 630014
rect 288942 629778 289026 630014
rect 289262 629778 289294 630014
rect 288674 596334 289294 629778
rect 288674 596098 288706 596334
rect 288942 596098 289026 596334
rect 289262 596098 289294 596334
rect 288674 596014 289294 596098
rect 288674 595778 288706 596014
rect 288942 595778 289026 596014
rect 289262 595778 289294 596014
rect 288674 562334 289294 595778
rect 288674 562098 288706 562334
rect 288942 562098 289026 562334
rect 289262 562098 289294 562334
rect 288674 562014 289294 562098
rect 288674 561778 288706 562014
rect 288942 561778 289026 562014
rect 289262 561778 289294 562014
rect 288674 528334 289294 561778
rect 288674 528098 288706 528334
rect 288942 528098 289026 528334
rect 289262 528098 289294 528334
rect 288674 528014 289294 528098
rect 288674 527778 288706 528014
rect 288942 527778 289026 528014
rect 289262 527778 289294 528014
rect 288674 494334 289294 527778
rect 288674 494098 288706 494334
rect 288942 494098 289026 494334
rect 289262 494098 289294 494334
rect 288674 494014 289294 494098
rect 288674 493778 288706 494014
rect 288942 493778 289026 494014
rect 289262 493778 289294 494014
rect 288674 460334 289294 493778
rect 288674 460098 288706 460334
rect 288942 460098 289026 460334
rect 289262 460098 289294 460334
rect 288674 460014 289294 460098
rect 288674 459778 288706 460014
rect 288942 459778 289026 460014
rect 289262 459778 289294 460014
rect 288674 426334 289294 459778
rect 288674 426098 288706 426334
rect 288942 426098 289026 426334
rect 289262 426098 289294 426334
rect 288674 426014 289294 426098
rect 288674 425778 288706 426014
rect 288942 425778 289026 426014
rect 289262 425778 289294 426014
rect 288674 392334 289294 425778
rect 288674 392098 288706 392334
rect 288942 392098 289026 392334
rect 289262 392098 289294 392334
rect 288674 392014 289294 392098
rect 288674 391778 288706 392014
rect 288942 391778 289026 392014
rect 289262 391778 289294 392014
rect 288674 358334 289294 391778
rect 288674 358098 288706 358334
rect 288942 358098 289026 358334
rect 289262 358098 289294 358334
rect 288674 358014 289294 358098
rect 288674 357778 288706 358014
rect 288942 357778 289026 358014
rect 289262 357778 289294 358014
rect 288674 324334 289294 357778
rect 288674 324098 288706 324334
rect 288942 324098 289026 324334
rect 289262 324098 289294 324334
rect 288674 324014 289294 324098
rect 288674 323778 288706 324014
rect 288942 323778 289026 324014
rect 289262 323778 289294 324014
rect 288674 290334 289294 323778
rect 288674 290098 288706 290334
rect 288942 290098 289026 290334
rect 289262 290098 289294 290334
rect 288674 290014 289294 290098
rect 288674 289778 288706 290014
rect 288942 289778 289026 290014
rect 289262 289778 289294 290014
rect 288674 256334 289294 289778
rect 288674 256098 288706 256334
rect 288942 256098 289026 256334
rect 289262 256098 289294 256334
rect 288674 256014 289294 256098
rect 288674 255778 288706 256014
rect 288942 255778 289026 256014
rect 289262 255778 289294 256014
rect 288674 225660 289294 255778
rect 292394 709638 293014 711590
rect 292394 709402 292426 709638
rect 292662 709402 292746 709638
rect 292982 709402 293014 709638
rect 292394 709318 293014 709402
rect 292394 709082 292426 709318
rect 292662 709082 292746 709318
rect 292982 709082 293014 709318
rect 292394 668054 293014 709082
rect 292394 667818 292426 668054
rect 292662 667818 292746 668054
rect 292982 667818 293014 668054
rect 292394 667734 293014 667818
rect 292394 667498 292426 667734
rect 292662 667498 292746 667734
rect 292982 667498 293014 667734
rect 292394 634054 293014 667498
rect 292394 633818 292426 634054
rect 292662 633818 292746 634054
rect 292982 633818 293014 634054
rect 292394 633734 293014 633818
rect 292394 633498 292426 633734
rect 292662 633498 292746 633734
rect 292982 633498 293014 633734
rect 292394 600054 293014 633498
rect 292394 599818 292426 600054
rect 292662 599818 292746 600054
rect 292982 599818 293014 600054
rect 292394 599734 293014 599818
rect 292394 599498 292426 599734
rect 292662 599498 292746 599734
rect 292982 599498 293014 599734
rect 292394 566054 293014 599498
rect 292394 565818 292426 566054
rect 292662 565818 292746 566054
rect 292982 565818 293014 566054
rect 292394 565734 293014 565818
rect 292394 565498 292426 565734
rect 292662 565498 292746 565734
rect 292982 565498 293014 565734
rect 292394 532054 293014 565498
rect 292394 531818 292426 532054
rect 292662 531818 292746 532054
rect 292982 531818 293014 532054
rect 292394 531734 293014 531818
rect 292394 531498 292426 531734
rect 292662 531498 292746 531734
rect 292982 531498 293014 531734
rect 292394 498054 293014 531498
rect 292394 497818 292426 498054
rect 292662 497818 292746 498054
rect 292982 497818 293014 498054
rect 292394 497734 293014 497818
rect 292394 497498 292426 497734
rect 292662 497498 292746 497734
rect 292982 497498 293014 497734
rect 292394 464054 293014 497498
rect 292394 463818 292426 464054
rect 292662 463818 292746 464054
rect 292982 463818 293014 464054
rect 292394 463734 293014 463818
rect 292394 463498 292426 463734
rect 292662 463498 292746 463734
rect 292982 463498 293014 463734
rect 292394 430054 293014 463498
rect 292394 429818 292426 430054
rect 292662 429818 292746 430054
rect 292982 429818 293014 430054
rect 292394 429734 293014 429818
rect 292394 429498 292426 429734
rect 292662 429498 292746 429734
rect 292982 429498 293014 429734
rect 292394 396054 293014 429498
rect 292394 395818 292426 396054
rect 292662 395818 292746 396054
rect 292982 395818 293014 396054
rect 292394 395734 293014 395818
rect 292394 395498 292426 395734
rect 292662 395498 292746 395734
rect 292982 395498 293014 395734
rect 292394 362054 293014 395498
rect 292394 361818 292426 362054
rect 292662 361818 292746 362054
rect 292982 361818 293014 362054
rect 292394 361734 293014 361818
rect 292394 361498 292426 361734
rect 292662 361498 292746 361734
rect 292982 361498 293014 361734
rect 292394 328054 293014 361498
rect 292394 327818 292426 328054
rect 292662 327818 292746 328054
rect 292982 327818 293014 328054
rect 292394 327734 293014 327818
rect 292394 327498 292426 327734
rect 292662 327498 292746 327734
rect 292982 327498 293014 327734
rect 292394 294054 293014 327498
rect 292394 293818 292426 294054
rect 292662 293818 292746 294054
rect 292982 293818 293014 294054
rect 292394 293734 293014 293818
rect 292394 293498 292426 293734
rect 292662 293498 292746 293734
rect 292982 293498 293014 293734
rect 292394 260054 293014 293498
rect 292394 259818 292426 260054
rect 292662 259818 292746 260054
rect 292982 259818 293014 260054
rect 292394 259734 293014 259818
rect 292394 259498 292426 259734
rect 292662 259498 292746 259734
rect 292982 259498 293014 259734
rect 292394 225991 293014 259498
rect 292394 225755 292426 225991
rect 292662 225755 292746 225991
rect 292982 225755 293014 225991
rect 292394 225660 293014 225755
rect 296114 710598 296734 711590
rect 296114 710362 296146 710598
rect 296382 710362 296466 710598
rect 296702 710362 296734 710598
rect 296114 710278 296734 710362
rect 296114 710042 296146 710278
rect 296382 710042 296466 710278
rect 296702 710042 296734 710278
rect 296114 671774 296734 710042
rect 296114 671538 296146 671774
rect 296382 671538 296466 671774
rect 296702 671538 296734 671774
rect 296114 671454 296734 671538
rect 296114 671218 296146 671454
rect 296382 671218 296466 671454
rect 296702 671218 296734 671454
rect 296114 637774 296734 671218
rect 296114 637538 296146 637774
rect 296382 637538 296466 637774
rect 296702 637538 296734 637774
rect 296114 637454 296734 637538
rect 296114 637218 296146 637454
rect 296382 637218 296466 637454
rect 296702 637218 296734 637454
rect 296114 603774 296734 637218
rect 296114 603538 296146 603774
rect 296382 603538 296466 603774
rect 296702 603538 296734 603774
rect 296114 603454 296734 603538
rect 296114 603218 296146 603454
rect 296382 603218 296466 603454
rect 296702 603218 296734 603454
rect 296114 569774 296734 603218
rect 296114 569538 296146 569774
rect 296382 569538 296466 569774
rect 296702 569538 296734 569774
rect 296114 569454 296734 569538
rect 296114 569218 296146 569454
rect 296382 569218 296466 569454
rect 296702 569218 296734 569454
rect 296114 535774 296734 569218
rect 296114 535538 296146 535774
rect 296382 535538 296466 535774
rect 296702 535538 296734 535774
rect 296114 535454 296734 535538
rect 296114 535218 296146 535454
rect 296382 535218 296466 535454
rect 296702 535218 296734 535454
rect 296114 501774 296734 535218
rect 296114 501538 296146 501774
rect 296382 501538 296466 501774
rect 296702 501538 296734 501774
rect 296114 501454 296734 501538
rect 296114 501218 296146 501454
rect 296382 501218 296466 501454
rect 296702 501218 296734 501454
rect 296114 467774 296734 501218
rect 296114 467538 296146 467774
rect 296382 467538 296466 467774
rect 296702 467538 296734 467774
rect 296114 467454 296734 467538
rect 296114 467218 296146 467454
rect 296382 467218 296466 467454
rect 296702 467218 296734 467454
rect 296114 433774 296734 467218
rect 296114 433538 296146 433774
rect 296382 433538 296466 433774
rect 296702 433538 296734 433774
rect 296114 433454 296734 433538
rect 296114 433218 296146 433454
rect 296382 433218 296466 433454
rect 296702 433218 296734 433454
rect 296114 399774 296734 433218
rect 296114 399538 296146 399774
rect 296382 399538 296466 399774
rect 296702 399538 296734 399774
rect 296114 399454 296734 399538
rect 296114 399218 296146 399454
rect 296382 399218 296466 399454
rect 296702 399218 296734 399454
rect 296114 365774 296734 399218
rect 296114 365538 296146 365774
rect 296382 365538 296466 365774
rect 296702 365538 296734 365774
rect 296114 365454 296734 365538
rect 296114 365218 296146 365454
rect 296382 365218 296466 365454
rect 296702 365218 296734 365454
rect 296114 331774 296734 365218
rect 296114 331538 296146 331774
rect 296382 331538 296466 331774
rect 296702 331538 296734 331774
rect 296114 331454 296734 331538
rect 296114 331218 296146 331454
rect 296382 331218 296466 331454
rect 296702 331218 296734 331454
rect 296114 297774 296734 331218
rect 296114 297538 296146 297774
rect 296382 297538 296466 297774
rect 296702 297538 296734 297774
rect 296114 297454 296734 297538
rect 296114 297218 296146 297454
rect 296382 297218 296466 297454
rect 296702 297218 296734 297454
rect 296114 263774 296734 297218
rect 296114 263538 296146 263774
rect 296382 263538 296466 263774
rect 296702 263538 296734 263774
rect 296114 263454 296734 263538
rect 296114 263218 296146 263454
rect 296382 263218 296466 263454
rect 296702 263218 296734 263454
rect 296114 229774 296734 263218
rect 296114 229538 296146 229774
rect 296382 229538 296466 229774
rect 296702 229538 296734 229774
rect 296114 229454 296734 229538
rect 296114 229218 296146 229454
rect 296382 229218 296466 229454
rect 296702 229218 296734 229454
rect 296114 225660 296734 229218
rect 299834 711558 300454 711590
rect 299834 711322 299866 711558
rect 300102 711322 300186 711558
rect 300422 711322 300454 711558
rect 299834 711238 300454 711322
rect 299834 711002 299866 711238
rect 300102 711002 300186 711238
rect 300422 711002 300454 711238
rect 299834 675494 300454 711002
rect 299834 675258 299866 675494
rect 300102 675258 300186 675494
rect 300422 675258 300454 675494
rect 299834 675174 300454 675258
rect 299834 674938 299866 675174
rect 300102 674938 300186 675174
rect 300422 674938 300454 675174
rect 299834 641494 300454 674938
rect 299834 641258 299866 641494
rect 300102 641258 300186 641494
rect 300422 641258 300454 641494
rect 299834 641174 300454 641258
rect 299834 640938 299866 641174
rect 300102 640938 300186 641174
rect 300422 640938 300454 641174
rect 299834 607494 300454 640938
rect 299834 607258 299866 607494
rect 300102 607258 300186 607494
rect 300422 607258 300454 607494
rect 299834 607174 300454 607258
rect 299834 606938 299866 607174
rect 300102 606938 300186 607174
rect 300422 606938 300454 607174
rect 299834 573494 300454 606938
rect 299834 573258 299866 573494
rect 300102 573258 300186 573494
rect 300422 573258 300454 573494
rect 299834 573174 300454 573258
rect 299834 572938 299866 573174
rect 300102 572938 300186 573174
rect 300422 572938 300454 573174
rect 299834 539494 300454 572938
rect 299834 539258 299866 539494
rect 300102 539258 300186 539494
rect 300422 539258 300454 539494
rect 299834 539174 300454 539258
rect 299834 538938 299866 539174
rect 300102 538938 300186 539174
rect 300422 538938 300454 539174
rect 299834 505494 300454 538938
rect 299834 505258 299866 505494
rect 300102 505258 300186 505494
rect 300422 505258 300454 505494
rect 299834 505174 300454 505258
rect 299834 504938 299866 505174
rect 300102 504938 300186 505174
rect 300422 504938 300454 505174
rect 299834 471494 300454 504938
rect 299834 471258 299866 471494
rect 300102 471258 300186 471494
rect 300422 471258 300454 471494
rect 299834 471174 300454 471258
rect 299834 470938 299866 471174
rect 300102 470938 300186 471174
rect 300422 470938 300454 471174
rect 299834 437494 300454 470938
rect 299834 437258 299866 437494
rect 300102 437258 300186 437494
rect 300422 437258 300454 437494
rect 299834 437174 300454 437258
rect 299834 436938 299866 437174
rect 300102 436938 300186 437174
rect 300422 436938 300454 437174
rect 299834 403494 300454 436938
rect 299834 403258 299866 403494
rect 300102 403258 300186 403494
rect 300422 403258 300454 403494
rect 299834 403174 300454 403258
rect 299834 402938 299866 403174
rect 300102 402938 300186 403174
rect 300422 402938 300454 403174
rect 299834 369494 300454 402938
rect 299834 369258 299866 369494
rect 300102 369258 300186 369494
rect 300422 369258 300454 369494
rect 299834 369174 300454 369258
rect 299834 368938 299866 369174
rect 300102 368938 300186 369174
rect 300422 368938 300454 369174
rect 299834 335494 300454 368938
rect 299834 335258 299866 335494
rect 300102 335258 300186 335494
rect 300422 335258 300454 335494
rect 299834 335174 300454 335258
rect 299834 334938 299866 335174
rect 300102 334938 300186 335174
rect 300422 334938 300454 335174
rect 299834 301494 300454 334938
rect 299834 301258 299866 301494
rect 300102 301258 300186 301494
rect 300422 301258 300454 301494
rect 299834 301174 300454 301258
rect 299834 300938 299866 301174
rect 300102 300938 300186 301174
rect 300422 300938 300454 301174
rect 299834 267494 300454 300938
rect 299834 267258 299866 267494
rect 300102 267258 300186 267494
rect 300422 267258 300454 267494
rect 299834 267174 300454 267258
rect 299834 266938 299866 267174
rect 300102 266938 300186 267174
rect 300422 266938 300454 267174
rect 299834 233494 300454 266938
rect 299834 233258 299866 233494
rect 300102 233258 300186 233494
rect 300422 233258 300454 233494
rect 299834 233174 300454 233258
rect 299834 232938 299866 233174
rect 300102 232938 300186 233174
rect 300422 232938 300454 233174
rect 299834 225660 300454 232938
rect 307794 704838 308414 711590
rect 307794 704602 307826 704838
rect 308062 704602 308146 704838
rect 308382 704602 308414 704838
rect 307794 704518 308414 704602
rect 307794 704282 307826 704518
rect 308062 704282 308146 704518
rect 308382 704282 308414 704518
rect 307794 683454 308414 704282
rect 307794 683218 307826 683454
rect 308062 683218 308146 683454
rect 308382 683218 308414 683454
rect 307794 683134 308414 683218
rect 307794 682898 307826 683134
rect 308062 682898 308146 683134
rect 308382 682898 308414 683134
rect 307794 649454 308414 682898
rect 307794 649218 307826 649454
rect 308062 649218 308146 649454
rect 308382 649218 308414 649454
rect 307794 649134 308414 649218
rect 307794 648898 307826 649134
rect 308062 648898 308146 649134
rect 308382 648898 308414 649134
rect 307794 615454 308414 648898
rect 307794 615218 307826 615454
rect 308062 615218 308146 615454
rect 308382 615218 308414 615454
rect 307794 615134 308414 615218
rect 307794 614898 307826 615134
rect 308062 614898 308146 615134
rect 308382 614898 308414 615134
rect 307794 581454 308414 614898
rect 307794 581218 307826 581454
rect 308062 581218 308146 581454
rect 308382 581218 308414 581454
rect 307794 581134 308414 581218
rect 307794 580898 307826 581134
rect 308062 580898 308146 581134
rect 308382 580898 308414 581134
rect 307794 547454 308414 580898
rect 307794 547218 307826 547454
rect 308062 547218 308146 547454
rect 308382 547218 308414 547454
rect 307794 547134 308414 547218
rect 307794 546898 307826 547134
rect 308062 546898 308146 547134
rect 308382 546898 308414 547134
rect 307794 513454 308414 546898
rect 307794 513218 307826 513454
rect 308062 513218 308146 513454
rect 308382 513218 308414 513454
rect 307794 513134 308414 513218
rect 307794 512898 307826 513134
rect 308062 512898 308146 513134
rect 308382 512898 308414 513134
rect 307794 479454 308414 512898
rect 307794 479218 307826 479454
rect 308062 479218 308146 479454
rect 308382 479218 308414 479454
rect 307794 479134 308414 479218
rect 307794 478898 307826 479134
rect 308062 478898 308146 479134
rect 308382 478898 308414 479134
rect 307794 445454 308414 478898
rect 307794 445218 307826 445454
rect 308062 445218 308146 445454
rect 308382 445218 308414 445454
rect 307794 445134 308414 445218
rect 307794 444898 307826 445134
rect 308062 444898 308146 445134
rect 308382 444898 308414 445134
rect 307794 411454 308414 444898
rect 307794 411218 307826 411454
rect 308062 411218 308146 411454
rect 308382 411218 308414 411454
rect 307794 411134 308414 411218
rect 307794 410898 307826 411134
rect 308062 410898 308146 411134
rect 308382 410898 308414 411134
rect 307794 377454 308414 410898
rect 307794 377218 307826 377454
rect 308062 377218 308146 377454
rect 308382 377218 308414 377454
rect 307794 377134 308414 377218
rect 307794 376898 307826 377134
rect 308062 376898 308146 377134
rect 308382 376898 308414 377134
rect 307794 343454 308414 376898
rect 307794 343218 307826 343454
rect 308062 343218 308146 343454
rect 308382 343218 308414 343454
rect 307794 343134 308414 343218
rect 307794 342898 307826 343134
rect 308062 342898 308146 343134
rect 308382 342898 308414 343134
rect 307794 309454 308414 342898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 275454 308414 308898
rect 307794 275218 307826 275454
rect 308062 275218 308146 275454
rect 308382 275218 308414 275454
rect 307794 275134 308414 275218
rect 307794 274898 307826 275134
rect 308062 274898 308146 275134
rect 308382 274898 308414 275134
rect 307794 241454 308414 274898
rect 307794 241218 307826 241454
rect 308062 241218 308146 241454
rect 308382 241218 308414 241454
rect 307794 241134 308414 241218
rect 307794 240898 307826 241134
rect 308062 240898 308146 241134
rect 308382 240898 308414 241134
rect 307794 225660 308414 240898
rect 311514 705798 312134 711590
rect 311514 705562 311546 705798
rect 311782 705562 311866 705798
rect 312102 705562 312134 705798
rect 311514 705478 312134 705562
rect 311514 705242 311546 705478
rect 311782 705242 311866 705478
rect 312102 705242 312134 705478
rect 311514 687174 312134 705242
rect 311514 686938 311546 687174
rect 311782 686938 311866 687174
rect 312102 686938 312134 687174
rect 311514 686854 312134 686938
rect 311514 686618 311546 686854
rect 311782 686618 311866 686854
rect 312102 686618 312134 686854
rect 311514 653174 312134 686618
rect 311514 652938 311546 653174
rect 311782 652938 311866 653174
rect 312102 652938 312134 653174
rect 311514 652854 312134 652938
rect 311514 652618 311546 652854
rect 311782 652618 311866 652854
rect 312102 652618 312134 652854
rect 311514 619174 312134 652618
rect 311514 618938 311546 619174
rect 311782 618938 311866 619174
rect 312102 618938 312134 619174
rect 311514 618854 312134 618938
rect 311514 618618 311546 618854
rect 311782 618618 311866 618854
rect 312102 618618 312134 618854
rect 311514 585174 312134 618618
rect 311514 584938 311546 585174
rect 311782 584938 311866 585174
rect 312102 584938 312134 585174
rect 311514 584854 312134 584938
rect 311514 584618 311546 584854
rect 311782 584618 311866 584854
rect 312102 584618 312134 584854
rect 311514 551174 312134 584618
rect 311514 550938 311546 551174
rect 311782 550938 311866 551174
rect 312102 550938 312134 551174
rect 311514 550854 312134 550938
rect 311514 550618 311546 550854
rect 311782 550618 311866 550854
rect 312102 550618 312134 550854
rect 311514 517174 312134 550618
rect 311514 516938 311546 517174
rect 311782 516938 311866 517174
rect 312102 516938 312134 517174
rect 311514 516854 312134 516938
rect 311514 516618 311546 516854
rect 311782 516618 311866 516854
rect 312102 516618 312134 516854
rect 311514 483174 312134 516618
rect 311514 482938 311546 483174
rect 311782 482938 311866 483174
rect 312102 482938 312134 483174
rect 311514 482854 312134 482938
rect 311514 482618 311546 482854
rect 311782 482618 311866 482854
rect 312102 482618 312134 482854
rect 311514 449174 312134 482618
rect 311514 448938 311546 449174
rect 311782 448938 311866 449174
rect 312102 448938 312134 449174
rect 311514 448854 312134 448938
rect 311514 448618 311546 448854
rect 311782 448618 311866 448854
rect 312102 448618 312134 448854
rect 311514 415174 312134 448618
rect 311514 414938 311546 415174
rect 311782 414938 311866 415174
rect 312102 414938 312134 415174
rect 311514 414854 312134 414938
rect 311514 414618 311546 414854
rect 311782 414618 311866 414854
rect 312102 414618 312134 414854
rect 311514 381174 312134 414618
rect 311514 380938 311546 381174
rect 311782 380938 311866 381174
rect 312102 380938 312134 381174
rect 311514 380854 312134 380938
rect 311514 380618 311546 380854
rect 311782 380618 311866 380854
rect 312102 380618 312134 380854
rect 311514 347174 312134 380618
rect 311514 346938 311546 347174
rect 311782 346938 311866 347174
rect 312102 346938 312134 347174
rect 311514 346854 312134 346938
rect 311514 346618 311546 346854
rect 311782 346618 311866 346854
rect 312102 346618 312134 346854
rect 311514 313174 312134 346618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 279174 312134 312618
rect 311514 278938 311546 279174
rect 311782 278938 311866 279174
rect 312102 278938 312134 279174
rect 311514 278854 312134 278938
rect 311514 278618 311546 278854
rect 311782 278618 311866 278854
rect 312102 278618 312134 278854
rect 311514 245174 312134 278618
rect 311514 244938 311546 245174
rect 311782 244938 311866 245174
rect 312102 244938 312134 245174
rect 311514 244854 312134 244938
rect 311514 244618 311546 244854
rect 311782 244618 311866 244854
rect 312102 244618 312134 244854
rect 281234 214658 281266 214894
rect 281502 214658 281586 214894
rect 281822 214658 281854 214894
rect 281234 214574 281854 214658
rect 250954 184378 250986 184614
rect 251222 184378 251306 184614
rect 251542 184378 251574 184614
rect 250954 184294 251574 184378
rect 250954 184058 250986 184294
rect 251222 184058 251306 184294
rect 251542 184058 251574 184294
rect 250954 150614 251574 184058
rect 250954 150378 250986 150614
rect 251222 150378 251306 150614
rect 251542 150378 251574 150614
rect 250954 150294 251574 150378
rect 250954 150058 250986 150294
rect 251222 150058 251306 150294
rect 251542 150058 251574 150294
rect 250954 116614 251574 150058
rect 250954 116378 250986 116614
rect 251222 116378 251306 116614
rect 251542 116378 251574 116614
rect 250954 116294 251574 116378
rect 250954 116058 250986 116294
rect 251222 116058 251306 116294
rect 251542 116058 251574 116294
rect 250954 82614 251574 116058
rect 250954 82378 250986 82614
rect 251222 82378 251306 82614
rect 251542 82378 251574 82614
rect 250954 82294 251574 82378
rect 250954 82058 250986 82294
rect 251222 82058 251306 82294
rect 251542 82058 251574 82294
rect 250954 48614 251574 82058
rect 250954 48378 250986 48614
rect 251222 48378 251306 48614
rect 251542 48378 251574 48614
rect 250954 48294 251574 48378
rect 250954 48058 250986 48294
rect 251222 48058 251306 48294
rect 251542 48058 251574 48294
rect 250954 14614 251574 48058
rect 250954 14378 250986 14614
rect 251222 14378 251306 14614
rect 251542 14378 251574 14614
rect 250954 14294 251574 14378
rect 250954 14058 250986 14294
rect 251222 14058 251306 14294
rect 251542 14058 251574 14294
rect 250954 -3226 251574 14058
rect 250954 -3462 250986 -3226
rect 251222 -3462 251306 -3226
rect 251542 -3462 251574 -3226
rect 250954 -3546 251574 -3462
rect 250954 -3782 250986 -3546
rect 251222 -3782 251306 -3546
rect 251542 -3782 251574 -3546
rect 250954 -7654 251574 -3782
rect 254674 188334 255294 214340
rect 254674 188098 254706 188334
rect 254942 188098 255026 188334
rect 255262 188098 255294 188334
rect 254674 188014 255294 188098
rect 254674 187778 254706 188014
rect 254942 187778 255026 188014
rect 255262 187778 255294 188014
rect 254674 154334 255294 187778
rect 254674 154098 254706 154334
rect 254942 154098 255026 154334
rect 255262 154098 255294 154334
rect 254674 154014 255294 154098
rect 254674 153778 254706 154014
rect 254942 153778 255026 154014
rect 255262 153778 255294 154014
rect 254674 120334 255294 153778
rect 254674 120098 254706 120334
rect 254942 120098 255026 120334
rect 255262 120098 255294 120334
rect 254674 120014 255294 120098
rect 254674 119778 254706 120014
rect 254942 119778 255026 120014
rect 255262 119778 255294 120014
rect 254674 86334 255294 119778
rect 254674 86098 254706 86334
rect 254942 86098 255026 86334
rect 255262 86098 255294 86334
rect 254674 86014 255294 86098
rect 254674 85778 254706 86014
rect 254942 85778 255026 86014
rect 255262 85778 255294 86014
rect 254674 52334 255294 85778
rect 254674 52098 254706 52334
rect 254942 52098 255026 52334
rect 255262 52098 255294 52334
rect 254674 52014 255294 52098
rect 254674 51778 254706 52014
rect 254942 51778 255026 52014
rect 255262 51778 255294 52014
rect 254674 18334 255294 51778
rect 254674 18098 254706 18334
rect 254942 18098 255026 18334
rect 255262 18098 255294 18334
rect 254674 18014 255294 18098
rect 254674 17778 254706 18014
rect 254942 17778 255026 18014
rect 255262 17778 255294 18014
rect 254674 -4186 255294 17778
rect 254674 -4422 254706 -4186
rect 254942 -4422 255026 -4186
rect 255262 -4422 255294 -4186
rect 254674 -4506 255294 -4422
rect 254674 -4742 254706 -4506
rect 254942 -4742 255026 -4506
rect 255262 -4742 255294 -4506
rect 254674 -7654 255294 -4742
rect 258394 192054 259014 214340
rect 258394 191818 258426 192054
rect 258662 191818 258746 192054
rect 258982 191818 259014 192054
rect 258394 191734 259014 191818
rect 258394 191498 258426 191734
rect 258662 191498 258746 191734
rect 258982 191498 259014 191734
rect 258394 158054 259014 191498
rect 258394 157818 258426 158054
rect 258662 157818 258746 158054
rect 258982 157818 259014 158054
rect 258394 157734 259014 157818
rect 258394 157498 258426 157734
rect 258662 157498 258746 157734
rect 258982 157498 259014 157734
rect 258394 124054 259014 157498
rect 258394 123818 258426 124054
rect 258662 123818 258746 124054
rect 258982 123818 259014 124054
rect 258394 123734 259014 123818
rect 258394 123498 258426 123734
rect 258662 123498 258746 123734
rect 258982 123498 259014 123734
rect 258394 90054 259014 123498
rect 258394 89818 258426 90054
rect 258662 89818 258746 90054
rect 258982 89818 259014 90054
rect 258394 89734 259014 89818
rect 258394 89498 258426 89734
rect 258662 89498 258746 89734
rect 258982 89498 259014 89734
rect 258394 56054 259014 89498
rect 258394 55818 258426 56054
rect 258662 55818 258746 56054
rect 258982 55818 259014 56054
rect 258394 55734 259014 55818
rect 258394 55498 258426 55734
rect 258662 55498 258746 55734
rect 258982 55498 259014 55734
rect 258394 22054 259014 55498
rect 258394 21818 258426 22054
rect 258662 21818 258746 22054
rect 258982 21818 259014 22054
rect 258394 21734 259014 21818
rect 258394 21498 258426 21734
rect 258662 21498 258746 21734
rect 258982 21498 259014 21734
rect 258394 -5146 259014 21498
rect 258394 -5382 258426 -5146
rect 258662 -5382 258746 -5146
rect 258982 -5382 259014 -5146
rect 258394 -5466 259014 -5382
rect 258394 -5702 258426 -5466
rect 258662 -5702 258746 -5466
rect 258982 -5702 259014 -5466
rect 258394 -7654 259014 -5702
rect 262114 195774 262734 214340
rect 262114 195538 262146 195774
rect 262382 195538 262466 195774
rect 262702 195538 262734 195774
rect 262114 195454 262734 195538
rect 262114 195218 262146 195454
rect 262382 195218 262466 195454
rect 262702 195218 262734 195454
rect 262114 161774 262734 195218
rect 262114 161538 262146 161774
rect 262382 161538 262466 161774
rect 262702 161538 262734 161774
rect 262114 161454 262734 161538
rect 262114 161218 262146 161454
rect 262382 161218 262466 161454
rect 262702 161218 262734 161454
rect 262114 127774 262734 161218
rect 262114 127538 262146 127774
rect 262382 127538 262466 127774
rect 262702 127538 262734 127774
rect 262114 127454 262734 127538
rect 262114 127218 262146 127454
rect 262382 127218 262466 127454
rect 262702 127218 262734 127454
rect 262114 93774 262734 127218
rect 262114 93538 262146 93774
rect 262382 93538 262466 93774
rect 262702 93538 262734 93774
rect 262114 93454 262734 93538
rect 262114 93218 262146 93454
rect 262382 93218 262466 93454
rect 262702 93218 262734 93454
rect 262114 59774 262734 93218
rect 262114 59538 262146 59774
rect 262382 59538 262466 59774
rect 262702 59538 262734 59774
rect 262114 59454 262734 59538
rect 262114 59218 262146 59454
rect 262382 59218 262466 59454
rect 262702 59218 262734 59454
rect 262114 25774 262734 59218
rect 262114 25538 262146 25774
rect 262382 25538 262466 25774
rect 262702 25538 262734 25774
rect 262114 25454 262734 25538
rect 262114 25218 262146 25454
rect 262382 25218 262466 25454
rect 262702 25218 262734 25454
rect 262114 -6106 262734 25218
rect 262114 -6342 262146 -6106
rect 262382 -6342 262466 -6106
rect 262702 -6342 262734 -6106
rect 262114 -6426 262734 -6342
rect 262114 -6662 262146 -6426
rect 262382 -6662 262466 -6426
rect 262702 -6662 262734 -6426
rect 262114 -7654 262734 -6662
rect 265834 199494 266454 214340
rect 265834 199258 265866 199494
rect 266102 199258 266186 199494
rect 266422 199258 266454 199494
rect 265834 199174 266454 199258
rect 265834 198938 265866 199174
rect 266102 198938 266186 199174
rect 266422 198938 266454 199174
rect 265834 165494 266454 198938
rect 265834 165258 265866 165494
rect 266102 165258 266186 165494
rect 266422 165258 266454 165494
rect 265834 165174 266454 165258
rect 265834 164938 265866 165174
rect 266102 164938 266186 165174
rect 266422 164938 266454 165174
rect 265834 131494 266454 164938
rect 265834 131258 265866 131494
rect 266102 131258 266186 131494
rect 266422 131258 266454 131494
rect 265834 131174 266454 131258
rect 265834 130938 265866 131174
rect 266102 130938 266186 131174
rect 266422 130938 266454 131174
rect 265834 97494 266454 130938
rect 265834 97258 265866 97494
rect 266102 97258 266186 97494
rect 266422 97258 266454 97494
rect 265834 97174 266454 97258
rect 265834 96938 265866 97174
rect 266102 96938 266186 97174
rect 266422 96938 266454 97174
rect 265834 63494 266454 96938
rect 265834 63258 265866 63494
rect 266102 63258 266186 63494
rect 266422 63258 266454 63494
rect 265834 63174 266454 63258
rect 265834 62938 265866 63174
rect 266102 62938 266186 63174
rect 266422 62938 266454 63174
rect 265834 29494 266454 62938
rect 265834 29258 265866 29494
rect 266102 29258 266186 29494
rect 266422 29258 266454 29494
rect 265834 29174 266454 29258
rect 265834 28938 265866 29174
rect 266102 28938 266186 29174
rect 266422 28938 266454 29174
rect 265834 -7066 266454 28938
rect 265834 -7302 265866 -7066
rect 266102 -7302 266186 -7066
rect 266422 -7302 266454 -7066
rect 265834 -7386 266454 -7302
rect 265834 -7622 265866 -7386
rect 266102 -7622 266186 -7386
rect 266422 -7622 266454 -7386
rect 265834 -7654 266454 -7622
rect 273794 207454 274414 214340
rect 273794 207218 273826 207454
rect 274062 207218 274146 207454
rect 274382 207218 274414 207454
rect 273794 207134 274414 207218
rect 273794 206898 273826 207134
rect 274062 206898 274146 207134
rect 274382 206898 274414 207134
rect 273794 173454 274414 206898
rect 273794 173218 273826 173454
rect 274062 173218 274146 173454
rect 274382 173218 274414 173454
rect 273794 173134 274414 173218
rect 273794 172898 273826 173134
rect 274062 172898 274146 173134
rect 274382 172898 274414 173134
rect 273794 139454 274414 172898
rect 273794 139218 273826 139454
rect 274062 139218 274146 139454
rect 274382 139218 274414 139454
rect 273794 139134 274414 139218
rect 273794 138898 273826 139134
rect 274062 138898 274146 139134
rect 274382 138898 274414 139134
rect 273794 105454 274414 138898
rect 273794 105218 273826 105454
rect 274062 105218 274146 105454
rect 274382 105218 274414 105454
rect 273794 105134 274414 105218
rect 273794 104898 273826 105134
rect 274062 104898 274146 105134
rect 274382 104898 274414 105134
rect 273794 71454 274414 104898
rect 273794 71218 273826 71454
rect 274062 71218 274146 71454
rect 274382 71218 274414 71454
rect 273794 71134 274414 71218
rect 273794 70898 273826 71134
rect 274062 70898 274146 71134
rect 274382 70898 274414 71134
rect 273794 37454 274414 70898
rect 273794 37218 273826 37454
rect 274062 37218 274146 37454
rect 274382 37218 274414 37454
rect 273794 37134 274414 37218
rect 273794 36898 273826 37134
rect 274062 36898 274146 37134
rect 274382 36898 274414 37134
rect 273794 3454 274414 36898
rect 273794 3218 273826 3454
rect 274062 3218 274146 3454
rect 274382 3218 274414 3454
rect 273794 3134 274414 3218
rect 273794 2898 273826 3134
rect 274062 2898 274146 3134
rect 274382 2898 274414 3134
rect 273794 -346 274414 2898
rect 273794 -582 273826 -346
rect 274062 -582 274146 -346
rect 274382 -582 274414 -346
rect 273794 -666 274414 -582
rect 273794 -902 273826 -666
rect 274062 -902 274146 -666
rect 274382 -902 274414 -666
rect 273794 -7654 274414 -902
rect 277514 211174 278134 214340
rect 277514 210938 277546 211174
rect 277782 210938 277866 211174
rect 278102 210938 278134 211174
rect 277514 210854 278134 210938
rect 277514 210618 277546 210854
rect 277782 210618 277866 210854
rect 278102 210618 278134 210854
rect 277514 177174 278134 210618
rect 277514 176938 277546 177174
rect 277782 176938 277866 177174
rect 278102 176938 278134 177174
rect 277514 176854 278134 176938
rect 277514 176618 277546 176854
rect 277782 176618 277866 176854
rect 278102 176618 278134 176854
rect 277514 143174 278134 176618
rect 277514 142938 277546 143174
rect 277782 142938 277866 143174
rect 278102 142938 278134 143174
rect 277514 142854 278134 142938
rect 277514 142618 277546 142854
rect 277782 142618 277866 142854
rect 278102 142618 278134 142854
rect 277514 109174 278134 142618
rect 277514 108938 277546 109174
rect 277782 108938 277866 109174
rect 278102 108938 278134 109174
rect 277514 108854 278134 108938
rect 277514 108618 277546 108854
rect 277782 108618 277866 108854
rect 278102 108618 278134 108854
rect 277514 75174 278134 108618
rect 277514 74938 277546 75174
rect 277782 74938 277866 75174
rect 278102 74938 278134 75174
rect 277514 74854 278134 74938
rect 277514 74618 277546 74854
rect 277782 74618 277866 74854
rect 278102 74618 278134 74854
rect 277514 41174 278134 74618
rect 277514 40938 277546 41174
rect 277782 40938 277866 41174
rect 278102 40938 278134 41174
rect 277514 40854 278134 40938
rect 277514 40618 277546 40854
rect 277782 40618 277866 40854
rect 278102 40618 278134 40854
rect 277514 7174 278134 40618
rect 277514 6938 277546 7174
rect 277782 6938 277866 7174
rect 278102 6938 278134 7174
rect 277514 6854 278134 6938
rect 277514 6618 277546 6854
rect 277782 6618 277866 6854
rect 278102 6618 278134 6854
rect 277514 -1306 278134 6618
rect 277514 -1542 277546 -1306
rect 277782 -1542 277866 -1306
rect 278102 -1542 278134 -1306
rect 277514 -1626 278134 -1542
rect 277514 -1862 277546 -1626
rect 277782 -1862 277866 -1626
rect 278102 -1862 278134 -1626
rect 277514 -7654 278134 -1862
rect 281234 214338 281266 214574
rect 281502 214338 281586 214574
rect 281822 214338 281854 214574
rect 281234 180894 281854 214338
rect 281234 180658 281266 180894
rect 281502 180658 281586 180894
rect 281822 180658 281854 180894
rect 281234 180574 281854 180658
rect 281234 180338 281266 180574
rect 281502 180338 281586 180574
rect 281822 180338 281854 180574
rect 281234 146894 281854 180338
rect 281234 146658 281266 146894
rect 281502 146658 281586 146894
rect 281822 146658 281854 146894
rect 281234 146574 281854 146658
rect 281234 146338 281266 146574
rect 281502 146338 281586 146574
rect 281822 146338 281854 146574
rect 281234 112894 281854 146338
rect 281234 112658 281266 112894
rect 281502 112658 281586 112894
rect 281822 112658 281854 112894
rect 281234 112574 281854 112658
rect 281234 112338 281266 112574
rect 281502 112338 281586 112574
rect 281822 112338 281854 112574
rect 281234 78894 281854 112338
rect 281234 78658 281266 78894
rect 281502 78658 281586 78894
rect 281822 78658 281854 78894
rect 281234 78574 281854 78658
rect 281234 78338 281266 78574
rect 281502 78338 281586 78574
rect 281822 78338 281854 78574
rect 281234 44894 281854 78338
rect 281234 44658 281266 44894
rect 281502 44658 281586 44894
rect 281822 44658 281854 44894
rect 281234 44574 281854 44658
rect 281234 44338 281266 44574
rect 281502 44338 281586 44574
rect 281822 44338 281854 44574
rect 281234 10894 281854 44338
rect 281234 10658 281266 10894
rect 281502 10658 281586 10894
rect 281822 10658 281854 10894
rect 281234 10574 281854 10658
rect 281234 10338 281266 10574
rect 281502 10338 281586 10574
rect 281822 10338 281854 10574
rect 281234 -2266 281854 10338
rect 281234 -2502 281266 -2266
rect 281502 -2502 281586 -2266
rect 281822 -2502 281854 -2266
rect 281234 -2586 281854 -2502
rect 281234 -2822 281266 -2586
rect 281502 -2822 281586 -2586
rect 281822 -2822 281854 -2586
rect 281234 -7654 281854 -2822
rect 284954 184614 285574 214340
rect 284954 184378 284986 184614
rect 285222 184378 285306 184614
rect 285542 184378 285574 184614
rect 284954 184294 285574 184378
rect 284954 184058 284986 184294
rect 285222 184058 285306 184294
rect 285542 184058 285574 184294
rect 284954 150614 285574 184058
rect 284954 150378 284986 150614
rect 285222 150378 285306 150614
rect 285542 150378 285574 150614
rect 284954 150294 285574 150378
rect 284954 150058 284986 150294
rect 285222 150058 285306 150294
rect 285542 150058 285574 150294
rect 284954 116614 285574 150058
rect 284954 116378 284986 116614
rect 285222 116378 285306 116614
rect 285542 116378 285574 116614
rect 284954 116294 285574 116378
rect 284954 116058 284986 116294
rect 285222 116058 285306 116294
rect 285542 116058 285574 116294
rect 284954 82614 285574 116058
rect 284954 82378 284986 82614
rect 285222 82378 285306 82614
rect 285542 82378 285574 82614
rect 284954 82294 285574 82378
rect 284954 82058 284986 82294
rect 285222 82058 285306 82294
rect 285542 82058 285574 82294
rect 284954 48614 285574 82058
rect 284954 48378 284986 48614
rect 285222 48378 285306 48614
rect 285542 48378 285574 48614
rect 284954 48294 285574 48378
rect 284954 48058 284986 48294
rect 285222 48058 285306 48294
rect 285542 48058 285574 48294
rect 284954 14614 285574 48058
rect 284954 14378 284986 14614
rect 285222 14378 285306 14614
rect 285542 14378 285574 14614
rect 284954 14294 285574 14378
rect 284954 14058 284986 14294
rect 285222 14058 285306 14294
rect 285542 14058 285574 14294
rect 284954 -3226 285574 14058
rect 284954 -3462 284986 -3226
rect 285222 -3462 285306 -3226
rect 285542 -3462 285574 -3226
rect 284954 -3546 285574 -3462
rect 284954 -3782 284986 -3546
rect 285222 -3782 285306 -3546
rect 285542 -3782 285574 -3546
rect 284954 -7654 285574 -3782
rect 288674 188334 289294 214340
rect 288674 188098 288706 188334
rect 288942 188098 289026 188334
rect 289262 188098 289294 188334
rect 288674 188014 289294 188098
rect 288674 187778 288706 188014
rect 288942 187778 289026 188014
rect 289262 187778 289294 188014
rect 288674 154334 289294 187778
rect 288674 154098 288706 154334
rect 288942 154098 289026 154334
rect 289262 154098 289294 154334
rect 288674 154014 289294 154098
rect 288674 153778 288706 154014
rect 288942 153778 289026 154014
rect 289262 153778 289294 154014
rect 288674 120334 289294 153778
rect 288674 120098 288706 120334
rect 288942 120098 289026 120334
rect 289262 120098 289294 120334
rect 288674 120014 289294 120098
rect 288674 119778 288706 120014
rect 288942 119778 289026 120014
rect 289262 119778 289294 120014
rect 288674 86334 289294 119778
rect 288674 86098 288706 86334
rect 288942 86098 289026 86334
rect 289262 86098 289294 86334
rect 288674 86014 289294 86098
rect 288674 85778 288706 86014
rect 288942 85778 289026 86014
rect 289262 85778 289294 86014
rect 288674 52334 289294 85778
rect 288674 52098 288706 52334
rect 288942 52098 289026 52334
rect 289262 52098 289294 52334
rect 288674 52014 289294 52098
rect 288674 51778 288706 52014
rect 288942 51778 289026 52014
rect 289262 51778 289294 52014
rect 288674 18334 289294 51778
rect 288674 18098 288706 18334
rect 288942 18098 289026 18334
rect 289262 18098 289294 18334
rect 288674 18014 289294 18098
rect 288674 17778 288706 18014
rect 288942 17778 289026 18014
rect 289262 17778 289294 18014
rect 288674 -4186 289294 17778
rect 288674 -4422 288706 -4186
rect 288942 -4422 289026 -4186
rect 289262 -4422 289294 -4186
rect 288674 -4506 289294 -4422
rect 288674 -4742 288706 -4506
rect 288942 -4742 289026 -4506
rect 289262 -4742 289294 -4506
rect 288674 -7654 289294 -4742
rect 292394 192054 293014 214340
rect 292394 191818 292426 192054
rect 292662 191818 292746 192054
rect 292982 191818 293014 192054
rect 292394 191734 293014 191818
rect 292394 191498 292426 191734
rect 292662 191498 292746 191734
rect 292982 191498 293014 191734
rect 292394 158054 293014 191498
rect 292394 157818 292426 158054
rect 292662 157818 292746 158054
rect 292982 157818 293014 158054
rect 292394 157734 293014 157818
rect 292394 157498 292426 157734
rect 292662 157498 292746 157734
rect 292982 157498 293014 157734
rect 292394 124054 293014 157498
rect 292394 123818 292426 124054
rect 292662 123818 292746 124054
rect 292982 123818 293014 124054
rect 292394 123734 293014 123818
rect 292394 123498 292426 123734
rect 292662 123498 292746 123734
rect 292982 123498 293014 123734
rect 292394 90054 293014 123498
rect 292394 89818 292426 90054
rect 292662 89818 292746 90054
rect 292982 89818 293014 90054
rect 292394 89734 293014 89818
rect 292394 89498 292426 89734
rect 292662 89498 292746 89734
rect 292982 89498 293014 89734
rect 292394 56054 293014 89498
rect 292394 55818 292426 56054
rect 292662 55818 292746 56054
rect 292982 55818 293014 56054
rect 292394 55734 293014 55818
rect 292394 55498 292426 55734
rect 292662 55498 292746 55734
rect 292982 55498 293014 55734
rect 292394 22054 293014 55498
rect 292394 21818 292426 22054
rect 292662 21818 292746 22054
rect 292982 21818 293014 22054
rect 292394 21734 293014 21818
rect 292394 21498 292426 21734
rect 292662 21498 292746 21734
rect 292982 21498 293014 21734
rect 292394 -5146 293014 21498
rect 292394 -5382 292426 -5146
rect 292662 -5382 292746 -5146
rect 292982 -5382 293014 -5146
rect 292394 -5466 293014 -5382
rect 292394 -5702 292426 -5466
rect 292662 -5702 292746 -5466
rect 292982 -5702 293014 -5466
rect 292394 -7654 293014 -5702
rect 296114 195774 296734 214340
rect 296114 195538 296146 195774
rect 296382 195538 296466 195774
rect 296702 195538 296734 195774
rect 296114 195454 296734 195538
rect 296114 195218 296146 195454
rect 296382 195218 296466 195454
rect 296702 195218 296734 195454
rect 296114 161774 296734 195218
rect 296114 161538 296146 161774
rect 296382 161538 296466 161774
rect 296702 161538 296734 161774
rect 296114 161454 296734 161538
rect 296114 161218 296146 161454
rect 296382 161218 296466 161454
rect 296702 161218 296734 161454
rect 296114 127774 296734 161218
rect 296114 127538 296146 127774
rect 296382 127538 296466 127774
rect 296702 127538 296734 127774
rect 296114 127454 296734 127538
rect 296114 127218 296146 127454
rect 296382 127218 296466 127454
rect 296702 127218 296734 127454
rect 296114 93774 296734 127218
rect 296114 93538 296146 93774
rect 296382 93538 296466 93774
rect 296702 93538 296734 93774
rect 296114 93454 296734 93538
rect 296114 93218 296146 93454
rect 296382 93218 296466 93454
rect 296702 93218 296734 93454
rect 296114 59774 296734 93218
rect 296114 59538 296146 59774
rect 296382 59538 296466 59774
rect 296702 59538 296734 59774
rect 296114 59454 296734 59538
rect 296114 59218 296146 59454
rect 296382 59218 296466 59454
rect 296702 59218 296734 59454
rect 296114 25774 296734 59218
rect 296114 25538 296146 25774
rect 296382 25538 296466 25774
rect 296702 25538 296734 25774
rect 296114 25454 296734 25538
rect 296114 25218 296146 25454
rect 296382 25218 296466 25454
rect 296702 25218 296734 25454
rect 296114 -6106 296734 25218
rect 296114 -6342 296146 -6106
rect 296382 -6342 296466 -6106
rect 296702 -6342 296734 -6106
rect 296114 -6426 296734 -6342
rect 296114 -6662 296146 -6426
rect 296382 -6662 296466 -6426
rect 296702 -6662 296734 -6426
rect 296114 -7654 296734 -6662
rect 299834 199494 300454 214340
rect 299834 199258 299866 199494
rect 300102 199258 300186 199494
rect 300422 199258 300454 199494
rect 299834 199174 300454 199258
rect 299834 198938 299866 199174
rect 300102 198938 300186 199174
rect 300422 198938 300454 199174
rect 299834 165494 300454 198938
rect 299834 165258 299866 165494
rect 300102 165258 300186 165494
rect 300422 165258 300454 165494
rect 299834 165174 300454 165258
rect 299834 164938 299866 165174
rect 300102 164938 300186 165174
rect 300422 164938 300454 165174
rect 299834 131494 300454 164938
rect 299834 131258 299866 131494
rect 300102 131258 300186 131494
rect 300422 131258 300454 131494
rect 299834 131174 300454 131258
rect 299834 130938 299866 131174
rect 300102 130938 300186 131174
rect 300422 130938 300454 131174
rect 299834 97494 300454 130938
rect 299834 97258 299866 97494
rect 300102 97258 300186 97494
rect 300422 97258 300454 97494
rect 299834 97174 300454 97258
rect 299834 96938 299866 97174
rect 300102 96938 300186 97174
rect 300422 96938 300454 97174
rect 299834 63494 300454 96938
rect 299834 63258 299866 63494
rect 300102 63258 300186 63494
rect 300422 63258 300454 63494
rect 299834 63174 300454 63258
rect 299834 62938 299866 63174
rect 300102 62938 300186 63174
rect 300422 62938 300454 63174
rect 299834 29494 300454 62938
rect 299834 29258 299866 29494
rect 300102 29258 300186 29494
rect 300422 29258 300454 29494
rect 299834 29174 300454 29258
rect 299834 28938 299866 29174
rect 300102 28938 300186 29174
rect 300422 28938 300454 29174
rect 299834 -7066 300454 28938
rect 299834 -7302 299866 -7066
rect 300102 -7302 300186 -7066
rect 300422 -7302 300454 -7066
rect 299834 -7386 300454 -7302
rect 299834 -7622 299866 -7386
rect 300102 -7622 300186 -7386
rect 300422 -7622 300454 -7386
rect 299834 -7654 300454 -7622
rect 307794 207454 308414 214340
rect 307794 207218 307826 207454
rect 308062 207218 308146 207454
rect 308382 207218 308414 207454
rect 307794 207134 308414 207218
rect 307794 206898 307826 207134
rect 308062 206898 308146 207134
rect 308382 206898 308414 207134
rect 307794 173454 308414 206898
rect 307794 173218 307826 173454
rect 308062 173218 308146 173454
rect 308382 173218 308414 173454
rect 307794 173134 308414 173218
rect 307794 172898 307826 173134
rect 308062 172898 308146 173134
rect 308382 172898 308414 173134
rect 307794 139454 308414 172898
rect 307794 139218 307826 139454
rect 308062 139218 308146 139454
rect 308382 139218 308414 139454
rect 307794 139134 308414 139218
rect 307794 138898 307826 139134
rect 308062 138898 308146 139134
rect 308382 138898 308414 139134
rect 307794 105454 308414 138898
rect 307794 105218 307826 105454
rect 308062 105218 308146 105454
rect 308382 105218 308414 105454
rect 307794 105134 308414 105218
rect 307794 104898 307826 105134
rect 308062 104898 308146 105134
rect 308382 104898 308414 105134
rect 307794 71454 308414 104898
rect 307794 71218 307826 71454
rect 308062 71218 308146 71454
rect 308382 71218 308414 71454
rect 307794 71134 308414 71218
rect 307794 70898 307826 71134
rect 308062 70898 308146 71134
rect 308382 70898 308414 71134
rect 307794 37454 308414 70898
rect 307794 37218 307826 37454
rect 308062 37218 308146 37454
rect 308382 37218 308414 37454
rect 307794 37134 308414 37218
rect 307794 36898 307826 37134
rect 308062 36898 308146 37134
rect 308382 36898 308414 37134
rect 307794 3454 308414 36898
rect 307794 3218 307826 3454
rect 308062 3218 308146 3454
rect 308382 3218 308414 3454
rect 307794 3134 308414 3218
rect 307794 2898 307826 3134
rect 308062 2898 308146 3134
rect 308382 2898 308414 3134
rect 307794 -346 308414 2898
rect 307794 -582 307826 -346
rect 308062 -582 308146 -346
rect 308382 -582 308414 -346
rect 307794 -666 308414 -582
rect 307794 -902 307826 -666
rect 308062 -902 308146 -666
rect 308382 -902 308414 -666
rect 307794 -7654 308414 -902
rect 311514 211174 312134 244618
rect 315234 706758 315854 711590
rect 315234 706522 315266 706758
rect 315502 706522 315586 706758
rect 315822 706522 315854 706758
rect 315234 706438 315854 706522
rect 315234 706202 315266 706438
rect 315502 706202 315586 706438
rect 315822 706202 315854 706438
rect 315234 690894 315854 706202
rect 315234 690658 315266 690894
rect 315502 690658 315586 690894
rect 315822 690658 315854 690894
rect 315234 690574 315854 690658
rect 315234 690338 315266 690574
rect 315502 690338 315586 690574
rect 315822 690338 315854 690574
rect 315234 656894 315854 690338
rect 315234 656658 315266 656894
rect 315502 656658 315586 656894
rect 315822 656658 315854 656894
rect 315234 656574 315854 656658
rect 315234 656338 315266 656574
rect 315502 656338 315586 656574
rect 315822 656338 315854 656574
rect 315234 622894 315854 656338
rect 315234 622658 315266 622894
rect 315502 622658 315586 622894
rect 315822 622658 315854 622894
rect 315234 622574 315854 622658
rect 315234 622338 315266 622574
rect 315502 622338 315586 622574
rect 315822 622338 315854 622574
rect 315234 588894 315854 622338
rect 315234 588658 315266 588894
rect 315502 588658 315586 588894
rect 315822 588658 315854 588894
rect 315234 588574 315854 588658
rect 315234 588338 315266 588574
rect 315502 588338 315586 588574
rect 315822 588338 315854 588574
rect 315234 554894 315854 588338
rect 315234 554658 315266 554894
rect 315502 554658 315586 554894
rect 315822 554658 315854 554894
rect 315234 554574 315854 554658
rect 315234 554338 315266 554574
rect 315502 554338 315586 554574
rect 315822 554338 315854 554574
rect 315234 520894 315854 554338
rect 315234 520658 315266 520894
rect 315502 520658 315586 520894
rect 315822 520658 315854 520894
rect 315234 520574 315854 520658
rect 315234 520338 315266 520574
rect 315502 520338 315586 520574
rect 315822 520338 315854 520574
rect 315234 486894 315854 520338
rect 315234 486658 315266 486894
rect 315502 486658 315586 486894
rect 315822 486658 315854 486894
rect 315234 486574 315854 486658
rect 315234 486338 315266 486574
rect 315502 486338 315586 486574
rect 315822 486338 315854 486574
rect 315234 452894 315854 486338
rect 315234 452658 315266 452894
rect 315502 452658 315586 452894
rect 315822 452658 315854 452894
rect 315234 452574 315854 452658
rect 315234 452338 315266 452574
rect 315502 452338 315586 452574
rect 315822 452338 315854 452574
rect 315234 418894 315854 452338
rect 315234 418658 315266 418894
rect 315502 418658 315586 418894
rect 315822 418658 315854 418894
rect 315234 418574 315854 418658
rect 315234 418338 315266 418574
rect 315502 418338 315586 418574
rect 315822 418338 315854 418574
rect 315234 384894 315854 418338
rect 315234 384658 315266 384894
rect 315502 384658 315586 384894
rect 315822 384658 315854 384894
rect 315234 384574 315854 384658
rect 315234 384338 315266 384574
rect 315502 384338 315586 384574
rect 315822 384338 315854 384574
rect 315234 350894 315854 384338
rect 315234 350658 315266 350894
rect 315502 350658 315586 350894
rect 315822 350658 315854 350894
rect 315234 350574 315854 350658
rect 315234 350338 315266 350574
rect 315502 350338 315586 350574
rect 315822 350338 315854 350574
rect 315234 316894 315854 350338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 282894 315854 316338
rect 315234 282658 315266 282894
rect 315502 282658 315586 282894
rect 315822 282658 315854 282894
rect 315234 282574 315854 282658
rect 315234 282338 315266 282574
rect 315502 282338 315586 282574
rect 315822 282338 315854 282574
rect 315234 248894 315854 282338
rect 315234 248658 315266 248894
rect 315502 248658 315586 248894
rect 315822 248658 315854 248894
rect 315234 248574 315854 248658
rect 315234 248338 315266 248574
rect 315502 248338 315586 248574
rect 315822 248338 315854 248574
rect 315234 225660 315854 248338
rect 318954 707718 319574 711590
rect 318954 707482 318986 707718
rect 319222 707482 319306 707718
rect 319542 707482 319574 707718
rect 318954 707398 319574 707482
rect 318954 707162 318986 707398
rect 319222 707162 319306 707398
rect 319542 707162 319574 707398
rect 318954 694614 319574 707162
rect 318954 694378 318986 694614
rect 319222 694378 319306 694614
rect 319542 694378 319574 694614
rect 318954 694294 319574 694378
rect 318954 694058 318986 694294
rect 319222 694058 319306 694294
rect 319542 694058 319574 694294
rect 318954 660614 319574 694058
rect 318954 660378 318986 660614
rect 319222 660378 319306 660614
rect 319542 660378 319574 660614
rect 318954 660294 319574 660378
rect 318954 660058 318986 660294
rect 319222 660058 319306 660294
rect 319542 660058 319574 660294
rect 318954 626614 319574 660058
rect 318954 626378 318986 626614
rect 319222 626378 319306 626614
rect 319542 626378 319574 626614
rect 318954 626294 319574 626378
rect 318954 626058 318986 626294
rect 319222 626058 319306 626294
rect 319542 626058 319574 626294
rect 318954 592614 319574 626058
rect 318954 592378 318986 592614
rect 319222 592378 319306 592614
rect 319542 592378 319574 592614
rect 318954 592294 319574 592378
rect 318954 592058 318986 592294
rect 319222 592058 319306 592294
rect 319542 592058 319574 592294
rect 318954 558614 319574 592058
rect 318954 558378 318986 558614
rect 319222 558378 319306 558614
rect 319542 558378 319574 558614
rect 318954 558294 319574 558378
rect 318954 558058 318986 558294
rect 319222 558058 319306 558294
rect 319542 558058 319574 558294
rect 318954 524614 319574 558058
rect 318954 524378 318986 524614
rect 319222 524378 319306 524614
rect 319542 524378 319574 524614
rect 318954 524294 319574 524378
rect 318954 524058 318986 524294
rect 319222 524058 319306 524294
rect 319542 524058 319574 524294
rect 318954 490614 319574 524058
rect 318954 490378 318986 490614
rect 319222 490378 319306 490614
rect 319542 490378 319574 490614
rect 318954 490294 319574 490378
rect 318954 490058 318986 490294
rect 319222 490058 319306 490294
rect 319542 490058 319574 490294
rect 318954 456614 319574 490058
rect 318954 456378 318986 456614
rect 319222 456378 319306 456614
rect 319542 456378 319574 456614
rect 318954 456294 319574 456378
rect 318954 456058 318986 456294
rect 319222 456058 319306 456294
rect 319542 456058 319574 456294
rect 318954 422614 319574 456058
rect 318954 422378 318986 422614
rect 319222 422378 319306 422614
rect 319542 422378 319574 422614
rect 318954 422294 319574 422378
rect 318954 422058 318986 422294
rect 319222 422058 319306 422294
rect 319542 422058 319574 422294
rect 318954 388614 319574 422058
rect 318954 388378 318986 388614
rect 319222 388378 319306 388614
rect 319542 388378 319574 388614
rect 318954 388294 319574 388378
rect 318954 388058 318986 388294
rect 319222 388058 319306 388294
rect 319542 388058 319574 388294
rect 318954 354614 319574 388058
rect 318954 354378 318986 354614
rect 319222 354378 319306 354614
rect 319542 354378 319574 354614
rect 318954 354294 319574 354378
rect 318954 354058 318986 354294
rect 319222 354058 319306 354294
rect 319542 354058 319574 354294
rect 318954 320614 319574 354058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 286614 319574 320058
rect 318954 286378 318986 286614
rect 319222 286378 319306 286614
rect 319542 286378 319574 286614
rect 318954 286294 319574 286378
rect 318954 286058 318986 286294
rect 319222 286058 319306 286294
rect 319542 286058 319574 286294
rect 318954 252614 319574 286058
rect 318954 252378 318986 252614
rect 319222 252378 319306 252614
rect 319542 252378 319574 252614
rect 318954 252294 319574 252378
rect 318954 252058 318986 252294
rect 319222 252058 319306 252294
rect 319542 252058 319574 252294
rect 318954 225660 319574 252058
rect 322674 708678 323294 711590
rect 322674 708442 322706 708678
rect 322942 708442 323026 708678
rect 323262 708442 323294 708678
rect 322674 708358 323294 708442
rect 322674 708122 322706 708358
rect 322942 708122 323026 708358
rect 323262 708122 323294 708358
rect 322674 698334 323294 708122
rect 322674 698098 322706 698334
rect 322942 698098 323026 698334
rect 323262 698098 323294 698334
rect 322674 698014 323294 698098
rect 322674 697778 322706 698014
rect 322942 697778 323026 698014
rect 323262 697778 323294 698014
rect 322674 664334 323294 697778
rect 322674 664098 322706 664334
rect 322942 664098 323026 664334
rect 323262 664098 323294 664334
rect 322674 664014 323294 664098
rect 322674 663778 322706 664014
rect 322942 663778 323026 664014
rect 323262 663778 323294 664014
rect 322674 630334 323294 663778
rect 322674 630098 322706 630334
rect 322942 630098 323026 630334
rect 323262 630098 323294 630334
rect 322674 630014 323294 630098
rect 322674 629778 322706 630014
rect 322942 629778 323026 630014
rect 323262 629778 323294 630014
rect 322674 596334 323294 629778
rect 322674 596098 322706 596334
rect 322942 596098 323026 596334
rect 323262 596098 323294 596334
rect 322674 596014 323294 596098
rect 322674 595778 322706 596014
rect 322942 595778 323026 596014
rect 323262 595778 323294 596014
rect 322674 562334 323294 595778
rect 322674 562098 322706 562334
rect 322942 562098 323026 562334
rect 323262 562098 323294 562334
rect 322674 562014 323294 562098
rect 322674 561778 322706 562014
rect 322942 561778 323026 562014
rect 323262 561778 323294 562014
rect 322674 528334 323294 561778
rect 322674 528098 322706 528334
rect 322942 528098 323026 528334
rect 323262 528098 323294 528334
rect 322674 528014 323294 528098
rect 322674 527778 322706 528014
rect 322942 527778 323026 528014
rect 323262 527778 323294 528014
rect 322674 494334 323294 527778
rect 322674 494098 322706 494334
rect 322942 494098 323026 494334
rect 323262 494098 323294 494334
rect 322674 494014 323294 494098
rect 322674 493778 322706 494014
rect 322942 493778 323026 494014
rect 323262 493778 323294 494014
rect 322674 460334 323294 493778
rect 322674 460098 322706 460334
rect 322942 460098 323026 460334
rect 323262 460098 323294 460334
rect 322674 460014 323294 460098
rect 322674 459778 322706 460014
rect 322942 459778 323026 460014
rect 323262 459778 323294 460014
rect 322674 426334 323294 459778
rect 322674 426098 322706 426334
rect 322942 426098 323026 426334
rect 323262 426098 323294 426334
rect 322674 426014 323294 426098
rect 322674 425778 322706 426014
rect 322942 425778 323026 426014
rect 323262 425778 323294 426014
rect 322674 392334 323294 425778
rect 322674 392098 322706 392334
rect 322942 392098 323026 392334
rect 323262 392098 323294 392334
rect 322674 392014 323294 392098
rect 322674 391778 322706 392014
rect 322942 391778 323026 392014
rect 323262 391778 323294 392014
rect 322674 358334 323294 391778
rect 322674 358098 322706 358334
rect 322942 358098 323026 358334
rect 323262 358098 323294 358334
rect 322674 358014 323294 358098
rect 322674 357778 322706 358014
rect 322942 357778 323026 358014
rect 323262 357778 323294 358014
rect 322674 324334 323294 357778
rect 322674 324098 322706 324334
rect 322942 324098 323026 324334
rect 323262 324098 323294 324334
rect 322674 324014 323294 324098
rect 322674 323778 322706 324014
rect 322942 323778 323026 324014
rect 323262 323778 323294 324014
rect 322674 290334 323294 323778
rect 322674 290098 322706 290334
rect 322942 290098 323026 290334
rect 323262 290098 323294 290334
rect 322674 290014 323294 290098
rect 322674 289778 322706 290014
rect 322942 289778 323026 290014
rect 323262 289778 323294 290014
rect 322674 256334 323294 289778
rect 322674 256098 322706 256334
rect 322942 256098 323026 256334
rect 323262 256098 323294 256334
rect 322674 256014 323294 256098
rect 322674 255778 322706 256014
rect 322942 255778 323026 256014
rect 323262 255778 323294 256014
rect 322674 225660 323294 255778
rect 326394 709638 327014 711590
rect 326394 709402 326426 709638
rect 326662 709402 326746 709638
rect 326982 709402 327014 709638
rect 326394 709318 327014 709402
rect 326394 709082 326426 709318
rect 326662 709082 326746 709318
rect 326982 709082 327014 709318
rect 326394 668054 327014 709082
rect 326394 667818 326426 668054
rect 326662 667818 326746 668054
rect 326982 667818 327014 668054
rect 326394 667734 327014 667818
rect 326394 667498 326426 667734
rect 326662 667498 326746 667734
rect 326982 667498 327014 667734
rect 326394 634054 327014 667498
rect 326394 633818 326426 634054
rect 326662 633818 326746 634054
rect 326982 633818 327014 634054
rect 326394 633734 327014 633818
rect 326394 633498 326426 633734
rect 326662 633498 326746 633734
rect 326982 633498 327014 633734
rect 326394 600054 327014 633498
rect 326394 599818 326426 600054
rect 326662 599818 326746 600054
rect 326982 599818 327014 600054
rect 326394 599734 327014 599818
rect 326394 599498 326426 599734
rect 326662 599498 326746 599734
rect 326982 599498 327014 599734
rect 326394 566054 327014 599498
rect 326394 565818 326426 566054
rect 326662 565818 326746 566054
rect 326982 565818 327014 566054
rect 326394 565734 327014 565818
rect 326394 565498 326426 565734
rect 326662 565498 326746 565734
rect 326982 565498 327014 565734
rect 326394 532054 327014 565498
rect 326394 531818 326426 532054
rect 326662 531818 326746 532054
rect 326982 531818 327014 532054
rect 326394 531734 327014 531818
rect 326394 531498 326426 531734
rect 326662 531498 326746 531734
rect 326982 531498 327014 531734
rect 326394 498054 327014 531498
rect 326394 497818 326426 498054
rect 326662 497818 326746 498054
rect 326982 497818 327014 498054
rect 326394 497734 327014 497818
rect 326394 497498 326426 497734
rect 326662 497498 326746 497734
rect 326982 497498 327014 497734
rect 326394 464054 327014 497498
rect 326394 463818 326426 464054
rect 326662 463818 326746 464054
rect 326982 463818 327014 464054
rect 326394 463734 327014 463818
rect 326394 463498 326426 463734
rect 326662 463498 326746 463734
rect 326982 463498 327014 463734
rect 326394 430054 327014 463498
rect 326394 429818 326426 430054
rect 326662 429818 326746 430054
rect 326982 429818 327014 430054
rect 326394 429734 327014 429818
rect 326394 429498 326426 429734
rect 326662 429498 326746 429734
rect 326982 429498 327014 429734
rect 326394 396054 327014 429498
rect 326394 395818 326426 396054
rect 326662 395818 326746 396054
rect 326982 395818 327014 396054
rect 326394 395734 327014 395818
rect 326394 395498 326426 395734
rect 326662 395498 326746 395734
rect 326982 395498 327014 395734
rect 326394 362054 327014 395498
rect 326394 361818 326426 362054
rect 326662 361818 326746 362054
rect 326982 361818 327014 362054
rect 326394 361734 327014 361818
rect 326394 361498 326426 361734
rect 326662 361498 326746 361734
rect 326982 361498 327014 361734
rect 326394 328054 327014 361498
rect 326394 327818 326426 328054
rect 326662 327818 326746 328054
rect 326982 327818 327014 328054
rect 326394 327734 327014 327818
rect 326394 327498 326426 327734
rect 326662 327498 326746 327734
rect 326982 327498 327014 327734
rect 326394 294054 327014 327498
rect 326394 293818 326426 294054
rect 326662 293818 326746 294054
rect 326982 293818 327014 294054
rect 326394 293734 327014 293818
rect 326394 293498 326426 293734
rect 326662 293498 326746 293734
rect 326982 293498 327014 293734
rect 326394 260054 327014 293498
rect 326394 259818 326426 260054
rect 326662 259818 326746 260054
rect 326982 259818 327014 260054
rect 326394 259734 327014 259818
rect 326394 259498 326426 259734
rect 326662 259498 326746 259734
rect 326982 259498 327014 259734
rect 326394 225991 327014 259498
rect 326394 225755 326426 225991
rect 326662 225755 326746 225991
rect 326982 225755 327014 225991
rect 326394 225660 327014 225755
rect 330114 710598 330734 711590
rect 330114 710362 330146 710598
rect 330382 710362 330466 710598
rect 330702 710362 330734 710598
rect 330114 710278 330734 710362
rect 330114 710042 330146 710278
rect 330382 710042 330466 710278
rect 330702 710042 330734 710278
rect 330114 671774 330734 710042
rect 330114 671538 330146 671774
rect 330382 671538 330466 671774
rect 330702 671538 330734 671774
rect 330114 671454 330734 671538
rect 330114 671218 330146 671454
rect 330382 671218 330466 671454
rect 330702 671218 330734 671454
rect 330114 637774 330734 671218
rect 330114 637538 330146 637774
rect 330382 637538 330466 637774
rect 330702 637538 330734 637774
rect 330114 637454 330734 637538
rect 330114 637218 330146 637454
rect 330382 637218 330466 637454
rect 330702 637218 330734 637454
rect 330114 603774 330734 637218
rect 330114 603538 330146 603774
rect 330382 603538 330466 603774
rect 330702 603538 330734 603774
rect 330114 603454 330734 603538
rect 330114 603218 330146 603454
rect 330382 603218 330466 603454
rect 330702 603218 330734 603454
rect 330114 569774 330734 603218
rect 330114 569538 330146 569774
rect 330382 569538 330466 569774
rect 330702 569538 330734 569774
rect 330114 569454 330734 569538
rect 330114 569218 330146 569454
rect 330382 569218 330466 569454
rect 330702 569218 330734 569454
rect 330114 535774 330734 569218
rect 330114 535538 330146 535774
rect 330382 535538 330466 535774
rect 330702 535538 330734 535774
rect 330114 535454 330734 535538
rect 330114 535218 330146 535454
rect 330382 535218 330466 535454
rect 330702 535218 330734 535454
rect 330114 501774 330734 535218
rect 330114 501538 330146 501774
rect 330382 501538 330466 501774
rect 330702 501538 330734 501774
rect 330114 501454 330734 501538
rect 330114 501218 330146 501454
rect 330382 501218 330466 501454
rect 330702 501218 330734 501454
rect 330114 467774 330734 501218
rect 330114 467538 330146 467774
rect 330382 467538 330466 467774
rect 330702 467538 330734 467774
rect 330114 467454 330734 467538
rect 330114 467218 330146 467454
rect 330382 467218 330466 467454
rect 330702 467218 330734 467454
rect 330114 433774 330734 467218
rect 330114 433538 330146 433774
rect 330382 433538 330466 433774
rect 330702 433538 330734 433774
rect 330114 433454 330734 433538
rect 330114 433218 330146 433454
rect 330382 433218 330466 433454
rect 330702 433218 330734 433454
rect 330114 399774 330734 433218
rect 330114 399538 330146 399774
rect 330382 399538 330466 399774
rect 330702 399538 330734 399774
rect 330114 399454 330734 399538
rect 330114 399218 330146 399454
rect 330382 399218 330466 399454
rect 330702 399218 330734 399454
rect 330114 365774 330734 399218
rect 330114 365538 330146 365774
rect 330382 365538 330466 365774
rect 330702 365538 330734 365774
rect 330114 365454 330734 365538
rect 330114 365218 330146 365454
rect 330382 365218 330466 365454
rect 330702 365218 330734 365454
rect 330114 331774 330734 365218
rect 330114 331538 330146 331774
rect 330382 331538 330466 331774
rect 330702 331538 330734 331774
rect 330114 331454 330734 331538
rect 330114 331218 330146 331454
rect 330382 331218 330466 331454
rect 330702 331218 330734 331454
rect 330114 297774 330734 331218
rect 330114 297538 330146 297774
rect 330382 297538 330466 297774
rect 330702 297538 330734 297774
rect 330114 297454 330734 297538
rect 330114 297218 330146 297454
rect 330382 297218 330466 297454
rect 330702 297218 330734 297454
rect 330114 263774 330734 297218
rect 330114 263538 330146 263774
rect 330382 263538 330466 263774
rect 330702 263538 330734 263774
rect 330114 263454 330734 263538
rect 330114 263218 330146 263454
rect 330382 263218 330466 263454
rect 330702 263218 330734 263454
rect 330114 229774 330734 263218
rect 330114 229538 330146 229774
rect 330382 229538 330466 229774
rect 330702 229538 330734 229774
rect 330114 229454 330734 229538
rect 330114 229218 330146 229454
rect 330382 229218 330466 229454
rect 330702 229218 330734 229454
rect 330114 225660 330734 229218
rect 333834 711558 334454 711590
rect 333834 711322 333866 711558
rect 334102 711322 334186 711558
rect 334422 711322 334454 711558
rect 333834 711238 334454 711322
rect 333834 711002 333866 711238
rect 334102 711002 334186 711238
rect 334422 711002 334454 711238
rect 333834 675494 334454 711002
rect 333834 675258 333866 675494
rect 334102 675258 334186 675494
rect 334422 675258 334454 675494
rect 333834 675174 334454 675258
rect 333834 674938 333866 675174
rect 334102 674938 334186 675174
rect 334422 674938 334454 675174
rect 333834 641494 334454 674938
rect 333834 641258 333866 641494
rect 334102 641258 334186 641494
rect 334422 641258 334454 641494
rect 333834 641174 334454 641258
rect 333834 640938 333866 641174
rect 334102 640938 334186 641174
rect 334422 640938 334454 641174
rect 333834 607494 334454 640938
rect 333834 607258 333866 607494
rect 334102 607258 334186 607494
rect 334422 607258 334454 607494
rect 333834 607174 334454 607258
rect 333834 606938 333866 607174
rect 334102 606938 334186 607174
rect 334422 606938 334454 607174
rect 333834 573494 334454 606938
rect 333834 573258 333866 573494
rect 334102 573258 334186 573494
rect 334422 573258 334454 573494
rect 333834 573174 334454 573258
rect 333834 572938 333866 573174
rect 334102 572938 334186 573174
rect 334422 572938 334454 573174
rect 333834 539494 334454 572938
rect 333834 539258 333866 539494
rect 334102 539258 334186 539494
rect 334422 539258 334454 539494
rect 333834 539174 334454 539258
rect 333834 538938 333866 539174
rect 334102 538938 334186 539174
rect 334422 538938 334454 539174
rect 333834 505494 334454 538938
rect 333834 505258 333866 505494
rect 334102 505258 334186 505494
rect 334422 505258 334454 505494
rect 333834 505174 334454 505258
rect 333834 504938 333866 505174
rect 334102 504938 334186 505174
rect 334422 504938 334454 505174
rect 333834 471494 334454 504938
rect 333834 471258 333866 471494
rect 334102 471258 334186 471494
rect 334422 471258 334454 471494
rect 333834 471174 334454 471258
rect 333834 470938 333866 471174
rect 334102 470938 334186 471174
rect 334422 470938 334454 471174
rect 333834 437494 334454 470938
rect 333834 437258 333866 437494
rect 334102 437258 334186 437494
rect 334422 437258 334454 437494
rect 333834 437174 334454 437258
rect 333834 436938 333866 437174
rect 334102 436938 334186 437174
rect 334422 436938 334454 437174
rect 333834 403494 334454 436938
rect 333834 403258 333866 403494
rect 334102 403258 334186 403494
rect 334422 403258 334454 403494
rect 333834 403174 334454 403258
rect 333834 402938 333866 403174
rect 334102 402938 334186 403174
rect 334422 402938 334454 403174
rect 333834 369494 334454 402938
rect 333834 369258 333866 369494
rect 334102 369258 334186 369494
rect 334422 369258 334454 369494
rect 333834 369174 334454 369258
rect 333834 368938 333866 369174
rect 334102 368938 334186 369174
rect 334422 368938 334454 369174
rect 333834 335494 334454 368938
rect 333834 335258 333866 335494
rect 334102 335258 334186 335494
rect 334422 335258 334454 335494
rect 333834 335174 334454 335258
rect 333834 334938 333866 335174
rect 334102 334938 334186 335174
rect 334422 334938 334454 335174
rect 333834 301494 334454 334938
rect 333834 301258 333866 301494
rect 334102 301258 334186 301494
rect 334422 301258 334454 301494
rect 333834 301174 334454 301258
rect 333834 300938 333866 301174
rect 334102 300938 334186 301174
rect 334422 300938 334454 301174
rect 333834 267494 334454 300938
rect 333834 267258 333866 267494
rect 334102 267258 334186 267494
rect 334422 267258 334454 267494
rect 333834 267174 334454 267258
rect 333834 266938 333866 267174
rect 334102 266938 334186 267174
rect 334422 266938 334454 267174
rect 333834 233494 334454 266938
rect 333834 233258 333866 233494
rect 334102 233258 334186 233494
rect 334422 233258 334454 233494
rect 333834 233174 334454 233258
rect 333834 232938 333866 233174
rect 334102 232938 334186 233174
rect 334422 232938 334454 233174
rect 333834 225660 334454 232938
rect 341794 704838 342414 711590
rect 341794 704602 341826 704838
rect 342062 704602 342146 704838
rect 342382 704602 342414 704838
rect 341794 704518 342414 704602
rect 341794 704282 341826 704518
rect 342062 704282 342146 704518
rect 342382 704282 342414 704518
rect 341794 683454 342414 704282
rect 341794 683218 341826 683454
rect 342062 683218 342146 683454
rect 342382 683218 342414 683454
rect 341794 683134 342414 683218
rect 341794 682898 341826 683134
rect 342062 682898 342146 683134
rect 342382 682898 342414 683134
rect 341794 649454 342414 682898
rect 341794 649218 341826 649454
rect 342062 649218 342146 649454
rect 342382 649218 342414 649454
rect 341794 649134 342414 649218
rect 341794 648898 341826 649134
rect 342062 648898 342146 649134
rect 342382 648898 342414 649134
rect 341794 615454 342414 648898
rect 341794 615218 341826 615454
rect 342062 615218 342146 615454
rect 342382 615218 342414 615454
rect 341794 615134 342414 615218
rect 341794 614898 341826 615134
rect 342062 614898 342146 615134
rect 342382 614898 342414 615134
rect 341794 581454 342414 614898
rect 341794 581218 341826 581454
rect 342062 581218 342146 581454
rect 342382 581218 342414 581454
rect 341794 581134 342414 581218
rect 341794 580898 341826 581134
rect 342062 580898 342146 581134
rect 342382 580898 342414 581134
rect 341794 547454 342414 580898
rect 341794 547218 341826 547454
rect 342062 547218 342146 547454
rect 342382 547218 342414 547454
rect 341794 547134 342414 547218
rect 341794 546898 341826 547134
rect 342062 546898 342146 547134
rect 342382 546898 342414 547134
rect 341794 513454 342414 546898
rect 341794 513218 341826 513454
rect 342062 513218 342146 513454
rect 342382 513218 342414 513454
rect 341794 513134 342414 513218
rect 341794 512898 341826 513134
rect 342062 512898 342146 513134
rect 342382 512898 342414 513134
rect 341794 479454 342414 512898
rect 341794 479218 341826 479454
rect 342062 479218 342146 479454
rect 342382 479218 342414 479454
rect 341794 479134 342414 479218
rect 341794 478898 341826 479134
rect 342062 478898 342146 479134
rect 342382 478898 342414 479134
rect 341794 445454 342414 478898
rect 341794 445218 341826 445454
rect 342062 445218 342146 445454
rect 342382 445218 342414 445454
rect 341794 445134 342414 445218
rect 341794 444898 341826 445134
rect 342062 444898 342146 445134
rect 342382 444898 342414 445134
rect 341794 411454 342414 444898
rect 341794 411218 341826 411454
rect 342062 411218 342146 411454
rect 342382 411218 342414 411454
rect 341794 411134 342414 411218
rect 341794 410898 341826 411134
rect 342062 410898 342146 411134
rect 342382 410898 342414 411134
rect 341794 377454 342414 410898
rect 341794 377218 341826 377454
rect 342062 377218 342146 377454
rect 342382 377218 342414 377454
rect 341794 377134 342414 377218
rect 341794 376898 341826 377134
rect 342062 376898 342146 377134
rect 342382 376898 342414 377134
rect 341794 343454 342414 376898
rect 341794 343218 341826 343454
rect 342062 343218 342146 343454
rect 342382 343218 342414 343454
rect 341794 343134 342414 343218
rect 341794 342898 341826 343134
rect 342062 342898 342146 343134
rect 342382 342898 342414 343134
rect 341794 309454 342414 342898
rect 341794 309218 341826 309454
rect 342062 309218 342146 309454
rect 342382 309218 342414 309454
rect 341794 309134 342414 309218
rect 341794 308898 341826 309134
rect 342062 308898 342146 309134
rect 342382 308898 342414 309134
rect 341794 275454 342414 308898
rect 341794 275218 341826 275454
rect 342062 275218 342146 275454
rect 342382 275218 342414 275454
rect 341794 275134 342414 275218
rect 341794 274898 341826 275134
rect 342062 274898 342146 275134
rect 342382 274898 342414 275134
rect 341794 241454 342414 274898
rect 341794 241218 341826 241454
rect 342062 241218 342146 241454
rect 342382 241218 342414 241454
rect 341794 241134 342414 241218
rect 341794 240898 341826 241134
rect 342062 240898 342146 241134
rect 342382 240898 342414 241134
rect 311514 210938 311546 211174
rect 311782 210938 311866 211174
rect 312102 210938 312134 211174
rect 311514 210854 312134 210938
rect 311514 210618 311546 210854
rect 311782 210618 311866 210854
rect 312102 210618 312134 210854
rect 311514 177174 312134 210618
rect 311514 176938 311546 177174
rect 311782 176938 311866 177174
rect 312102 176938 312134 177174
rect 311514 176854 312134 176938
rect 311514 176618 311546 176854
rect 311782 176618 311866 176854
rect 312102 176618 312134 176854
rect 311514 143174 312134 176618
rect 311514 142938 311546 143174
rect 311782 142938 311866 143174
rect 312102 142938 312134 143174
rect 311514 142854 312134 142938
rect 311514 142618 311546 142854
rect 311782 142618 311866 142854
rect 312102 142618 312134 142854
rect 311514 109174 312134 142618
rect 311514 108938 311546 109174
rect 311782 108938 311866 109174
rect 312102 108938 312134 109174
rect 311514 108854 312134 108938
rect 311514 108618 311546 108854
rect 311782 108618 311866 108854
rect 312102 108618 312134 108854
rect 311514 75174 312134 108618
rect 311514 74938 311546 75174
rect 311782 74938 311866 75174
rect 312102 74938 312134 75174
rect 311514 74854 312134 74938
rect 311514 74618 311546 74854
rect 311782 74618 311866 74854
rect 312102 74618 312134 74854
rect 311514 41174 312134 74618
rect 311514 40938 311546 41174
rect 311782 40938 311866 41174
rect 312102 40938 312134 41174
rect 311514 40854 312134 40938
rect 311514 40618 311546 40854
rect 311782 40618 311866 40854
rect 312102 40618 312134 40854
rect 311514 7174 312134 40618
rect 311514 6938 311546 7174
rect 311782 6938 311866 7174
rect 312102 6938 312134 7174
rect 311514 6854 312134 6938
rect 311514 6618 311546 6854
rect 311782 6618 311866 6854
rect 312102 6618 312134 6854
rect 311514 -1306 312134 6618
rect 311514 -1542 311546 -1306
rect 311782 -1542 311866 -1306
rect 312102 -1542 312134 -1306
rect 311514 -1626 312134 -1542
rect 311514 -1862 311546 -1626
rect 311782 -1862 311866 -1626
rect 312102 -1862 312134 -1626
rect 311514 -7654 312134 -1862
rect 315234 180894 315854 214340
rect 315234 180658 315266 180894
rect 315502 180658 315586 180894
rect 315822 180658 315854 180894
rect 315234 180574 315854 180658
rect 315234 180338 315266 180574
rect 315502 180338 315586 180574
rect 315822 180338 315854 180574
rect 315234 146894 315854 180338
rect 315234 146658 315266 146894
rect 315502 146658 315586 146894
rect 315822 146658 315854 146894
rect 315234 146574 315854 146658
rect 315234 146338 315266 146574
rect 315502 146338 315586 146574
rect 315822 146338 315854 146574
rect 315234 112894 315854 146338
rect 315234 112658 315266 112894
rect 315502 112658 315586 112894
rect 315822 112658 315854 112894
rect 315234 112574 315854 112658
rect 315234 112338 315266 112574
rect 315502 112338 315586 112574
rect 315822 112338 315854 112574
rect 315234 78894 315854 112338
rect 315234 78658 315266 78894
rect 315502 78658 315586 78894
rect 315822 78658 315854 78894
rect 315234 78574 315854 78658
rect 315234 78338 315266 78574
rect 315502 78338 315586 78574
rect 315822 78338 315854 78574
rect 315234 44894 315854 78338
rect 315234 44658 315266 44894
rect 315502 44658 315586 44894
rect 315822 44658 315854 44894
rect 315234 44574 315854 44658
rect 315234 44338 315266 44574
rect 315502 44338 315586 44574
rect 315822 44338 315854 44574
rect 315234 10894 315854 44338
rect 315234 10658 315266 10894
rect 315502 10658 315586 10894
rect 315822 10658 315854 10894
rect 315234 10574 315854 10658
rect 315234 10338 315266 10574
rect 315502 10338 315586 10574
rect 315822 10338 315854 10574
rect 315234 -2266 315854 10338
rect 315234 -2502 315266 -2266
rect 315502 -2502 315586 -2266
rect 315822 -2502 315854 -2266
rect 315234 -2586 315854 -2502
rect 315234 -2822 315266 -2586
rect 315502 -2822 315586 -2586
rect 315822 -2822 315854 -2586
rect 315234 -7654 315854 -2822
rect 318954 184614 319574 214340
rect 318954 184378 318986 184614
rect 319222 184378 319306 184614
rect 319542 184378 319574 184614
rect 318954 184294 319574 184378
rect 318954 184058 318986 184294
rect 319222 184058 319306 184294
rect 319542 184058 319574 184294
rect 318954 150614 319574 184058
rect 318954 150378 318986 150614
rect 319222 150378 319306 150614
rect 319542 150378 319574 150614
rect 318954 150294 319574 150378
rect 318954 150058 318986 150294
rect 319222 150058 319306 150294
rect 319542 150058 319574 150294
rect 318954 116614 319574 150058
rect 318954 116378 318986 116614
rect 319222 116378 319306 116614
rect 319542 116378 319574 116614
rect 318954 116294 319574 116378
rect 318954 116058 318986 116294
rect 319222 116058 319306 116294
rect 319542 116058 319574 116294
rect 318954 82614 319574 116058
rect 318954 82378 318986 82614
rect 319222 82378 319306 82614
rect 319542 82378 319574 82614
rect 318954 82294 319574 82378
rect 318954 82058 318986 82294
rect 319222 82058 319306 82294
rect 319542 82058 319574 82294
rect 318954 48614 319574 82058
rect 318954 48378 318986 48614
rect 319222 48378 319306 48614
rect 319542 48378 319574 48614
rect 318954 48294 319574 48378
rect 318954 48058 318986 48294
rect 319222 48058 319306 48294
rect 319542 48058 319574 48294
rect 318954 14614 319574 48058
rect 318954 14378 318986 14614
rect 319222 14378 319306 14614
rect 319542 14378 319574 14614
rect 318954 14294 319574 14378
rect 318954 14058 318986 14294
rect 319222 14058 319306 14294
rect 319542 14058 319574 14294
rect 318954 -3226 319574 14058
rect 318954 -3462 318986 -3226
rect 319222 -3462 319306 -3226
rect 319542 -3462 319574 -3226
rect 318954 -3546 319574 -3462
rect 318954 -3782 318986 -3546
rect 319222 -3782 319306 -3546
rect 319542 -3782 319574 -3546
rect 318954 -7654 319574 -3782
rect 322674 188334 323294 214340
rect 322674 188098 322706 188334
rect 322942 188098 323026 188334
rect 323262 188098 323294 188334
rect 322674 188014 323294 188098
rect 322674 187778 322706 188014
rect 322942 187778 323026 188014
rect 323262 187778 323294 188014
rect 322674 154334 323294 187778
rect 322674 154098 322706 154334
rect 322942 154098 323026 154334
rect 323262 154098 323294 154334
rect 322674 154014 323294 154098
rect 322674 153778 322706 154014
rect 322942 153778 323026 154014
rect 323262 153778 323294 154014
rect 322674 120334 323294 153778
rect 322674 120098 322706 120334
rect 322942 120098 323026 120334
rect 323262 120098 323294 120334
rect 322674 120014 323294 120098
rect 322674 119778 322706 120014
rect 322942 119778 323026 120014
rect 323262 119778 323294 120014
rect 322674 86334 323294 119778
rect 322674 86098 322706 86334
rect 322942 86098 323026 86334
rect 323262 86098 323294 86334
rect 322674 86014 323294 86098
rect 322674 85778 322706 86014
rect 322942 85778 323026 86014
rect 323262 85778 323294 86014
rect 322674 52334 323294 85778
rect 322674 52098 322706 52334
rect 322942 52098 323026 52334
rect 323262 52098 323294 52334
rect 322674 52014 323294 52098
rect 322674 51778 322706 52014
rect 322942 51778 323026 52014
rect 323262 51778 323294 52014
rect 322674 18334 323294 51778
rect 322674 18098 322706 18334
rect 322942 18098 323026 18334
rect 323262 18098 323294 18334
rect 322674 18014 323294 18098
rect 322674 17778 322706 18014
rect 322942 17778 323026 18014
rect 323262 17778 323294 18014
rect 322674 -4186 323294 17778
rect 322674 -4422 322706 -4186
rect 322942 -4422 323026 -4186
rect 323262 -4422 323294 -4186
rect 322674 -4506 323294 -4422
rect 322674 -4742 322706 -4506
rect 322942 -4742 323026 -4506
rect 323262 -4742 323294 -4506
rect 322674 -7654 323294 -4742
rect 326394 192054 327014 214340
rect 326394 191818 326426 192054
rect 326662 191818 326746 192054
rect 326982 191818 327014 192054
rect 326394 191734 327014 191818
rect 326394 191498 326426 191734
rect 326662 191498 326746 191734
rect 326982 191498 327014 191734
rect 326394 158054 327014 191498
rect 326394 157818 326426 158054
rect 326662 157818 326746 158054
rect 326982 157818 327014 158054
rect 326394 157734 327014 157818
rect 326394 157498 326426 157734
rect 326662 157498 326746 157734
rect 326982 157498 327014 157734
rect 326394 124054 327014 157498
rect 326394 123818 326426 124054
rect 326662 123818 326746 124054
rect 326982 123818 327014 124054
rect 326394 123734 327014 123818
rect 326394 123498 326426 123734
rect 326662 123498 326746 123734
rect 326982 123498 327014 123734
rect 326394 90054 327014 123498
rect 326394 89818 326426 90054
rect 326662 89818 326746 90054
rect 326982 89818 327014 90054
rect 326394 89734 327014 89818
rect 326394 89498 326426 89734
rect 326662 89498 326746 89734
rect 326982 89498 327014 89734
rect 326394 56054 327014 89498
rect 326394 55818 326426 56054
rect 326662 55818 326746 56054
rect 326982 55818 327014 56054
rect 326394 55734 327014 55818
rect 326394 55498 326426 55734
rect 326662 55498 326746 55734
rect 326982 55498 327014 55734
rect 326394 22054 327014 55498
rect 326394 21818 326426 22054
rect 326662 21818 326746 22054
rect 326982 21818 327014 22054
rect 326394 21734 327014 21818
rect 326394 21498 326426 21734
rect 326662 21498 326746 21734
rect 326982 21498 327014 21734
rect 326394 -5146 327014 21498
rect 326394 -5382 326426 -5146
rect 326662 -5382 326746 -5146
rect 326982 -5382 327014 -5146
rect 326394 -5466 327014 -5382
rect 326394 -5702 326426 -5466
rect 326662 -5702 326746 -5466
rect 326982 -5702 327014 -5466
rect 326394 -7654 327014 -5702
rect 330114 195774 330734 214340
rect 330114 195538 330146 195774
rect 330382 195538 330466 195774
rect 330702 195538 330734 195774
rect 330114 195454 330734 195538
rect 330114 195218 330146 195454
rect 330382 195218 330466 195454
rect 330702 195218 330734 195454
rect 330114 161774 330734 195218
rect 330114 161538 330146 161774
rect 330382 161538 330466 161774
rect 330702 161538 330734 161774
rect 330114 161454 330734 161538
rect 330114 161218 330146 161454
rect 330382 161218 330466 161454
rect 330702 161218 330734 161454
rect 330114 127774 330734 161218
rect 330114 127538 330146 127774
rect 330382 127538 330466 127774
rect 330702 127538 330734 127774
rect 330114 127454 330734 127538
rect 330114 127218 330146 127454
rect 330382 127218 330466 127454
rect 330702 127218 330734 127454
rect 330114 93774 330734 127218
rect 330114 93538 330146 93774
rect 330382 93538 330466 93774
rect 330702 93538 330734 93774
rect 330114 93454 330734 93538
rect 330114 93218 330146 93454
rect 330382 93218 330466 93454
rect 330702 93218 330734 93454
rect 330114 59774 330734 93218
rect 330114 59538 330146 59774
rect 330382 59538 330466 59774
rect 330702 59538 330734 59774
rect 330114 59454 330734 59538
rect 330114 59218 330146 59454
rect 330382 59218 330466 59454
rect 330702 59218 330734 59454
rect 330114 25774 330734 59218
rect 330114 25538 330146 25774
rect 330382 25538 330466 25774
rect 330702 25538 330734 25774
rect 330114 25454 330734 25538
rect 330114 25218 330146 25454
rect 330382 25218 330466 25454
rect 330702 25218 330734 25454
rect 330114 -6106 330734 25218
rect 330114 -6342 330146 -6106
rect 330382 -6342 330466 -6106
rect 330702 -6342 330734 -6106
rect 330114 -6426 330734 -6342
rect 330114 -6662 330146 -6426
rect 330382 -6662 330466 -6426
rect 330702 -6662 330734 -6426
rect 330114 -7654 330734 -6662
rect 333834 199494 334454 214340
rect 333834 199258 333866 199494
rect 334102 199258 334186 199494
rect 334422 199258 334454 199494
rect 333834 199174 334454 199258
rect 333834 198938 333866 199174
rect 334102 198938 334186 199174
rect 334422 198938 334454 199174
rect 333834 165494 334454 198938
rect 333834 165258 333866 165494
rect 334102 165258 334186 165494
rect 334422 165258 334454 165494
rect 333834 165174 334454 165258
rect 333834 164938 333866 165174
rect 334102 164938 334186 165174
rect 334422 164938 334454 165174
rect 333834 131494 334454 164938
rect 333834 131258 333866 131494
rect 334102 131258 334186 131494
rect 334422 131258 334454 131494
rect 333834 131174 334454 131258
rect 333834 130938 333866 131174
rect 334102 130938 334186 131174
rect 334422 130938 334454 131174
rect 333834 97494 334454 130938
rect 333834 97258 333866 97494
rect 334102 97258 334186 97494
rect 334422 97258 334454 97494
rect 333834 97174 334454 97258
rect 333834 96938 333866 97174
rect 334102 96938 334186 97174
rect 334422 96938 334454 97174
rect 333834 63494 334454 96938
rect 333834 63258 333866 63494
rect 334102 63258 334186 63494
rect 334422 63258 334454 63494
rect 333834 63174 334454 63258
rect 333834 62938 333866 63174
rect 334102 62938 334186 63174
rect 334422 62938 334454 63174
rect 333834 29494 334454 62938
rect 333834 29258 333866 29494
rect 334102 29258 334186 29494
rect 334422 29258 334454 29494
rect 333834 29174 334454 29258
rect 333834 28938 333866 29174
rect 334102 28938 334186 29174
rect 334422 28938 334454 29174
rect 333834 -7066 334454 28938
rect 333834 -7302 333866 -7066
rect 334102 -7302 334186 -7066
rect 334422 -7302 334454 -7066
rect 333834 -7386 334454 -7302
rect 333834 -7622 333866 -7386
rect 334102 -7622 334186 -7386
rect 334422 -7622 334454 -7386
rect 333834 -7654 334454 -7622
rect 341794 207454 342414 240898
rect 345514 705798 346134 711590
rect 345514 705562 345546 705798
rect 345782 705562 345866 705798
rect 346102 705562 346134 705798
rect 345514 705478 346134 705562
rect 345514 705242 345546 705478
rect 345782 705242 345866 705478
rect 346102 705242 346134 705478
rect 345514 687174 346134 705242
rect 345514 686938 345546 687174
rect 345782 686938 345866 687174
rect 346102 686938 346134 687174
rect 345514 686854 346134 686938
rect 345514 686618 345546 686854
rect 345782 686618 345866 686854
rect 346102 686618 346134 686854
rect 345514 653174 346134 686618
rect 345514 652938 345546 653174
rect 345782 652938 345866 653174
rect 346102 652938 346134 653174
rect 345514 652854 346134 652938
rect 345514 652618 345546 652854
rect 345782 652618 345866 652854
rect 346102 652618 346134 652854
rect 345514 619174 346134 652618
rect 345514 618938 345546 619174
rect 345782 618938 345866 619174
rect 346102 618938 346134 619174
rect 345514 618854 346134 618938
rect 345514 618618 345546 618854
rect 345782 618618 345866 618854
rect 346102 618618 346134 618854
rect 345514 585174 346134 618618
rect 345514 584938 345546 585174
rect 345782 584938 345866 585174
rect 346102 584938 346134 585174
rect 345514 584854 346134 584938
rect 345514 584618 345546 584854
rect 345782 584618 345866 584854
rect 346102 584618 346134 584854
rect 345514 551174 346134 584618
rect 345514 550938 345546 551174
rect 345782 550938 345866 551174
rect 346102 550938 346134 551174
rect 345514 550854 346134 550938
rect 345514 550618 345546 550854
rect 345782 550618 345866 550854
rect 346102 550618 346134 550854
rect 345514 517174 346134 550618
rect 345514 516938 345546 517174
rect 345782 516938 345866 517174
rect 346102 516938 346134 517174
rect 345514 516854 346134 516938
rect 345514 516618 345546 516854
rect 345782 516618 345866 516854
rect 346102 516618 346134 516854
rect 345514 483174 346134 516618
rect 345514 482938 345546 483174
rect 345782 482938 345866 483174
rect 346102 482938 346134 483174
rect 345514 482854 346134 482938
rect 345514 482618 345546 482854
rect 345782 482618 345866 482854
rect 346102 482618 346134 482854
rect 345514 449174 346134 482618
rect 345514 448938 345546 449174
rect 345782 448938 345866 449174
rect 346102 448938 346134 449174
rect 345514 448854 346134 448938
rect 345514 448618 345546 448854
rect 345782 448618 345866 448854
rect 346102 448618 346134 448854
rect 345514 415174 346134 448618
rect 345514 414938 345546 415174
rect 345782 414938 345866 415174
rect 346102 414938 346134 415174
rect 345514 414854 346134 414938
rect 345514 414618 345546 414854
rect 345782 414618 345866 414854
rect 346102 414618 346134 414854
rect 345514 381174 346134 414618
rect 345514 380938 345546 381174
rect 345782 380938 345866 381174
rect 346102 380938 346134 381174
rect 345514 380854 346134 380938
rect 345514 380618 345546 380854
rect 345782 380618 345866 380854
rect 346102 380618 346134 380854
rect 345514 347174 346134 380618
rect 345514 346938 345546 347174
rect 345782 346938 345866 347174
rect 346102 346938 346134 347174
rect 345514 346854 346134 346938
rect 345514 346618 345546 346854
rect 345782 346618 345866 346854
rect 346102 346618 346134 346854
rect 345514 313174 346134 346618
rect 345514 312938 345546 313174
rect 345782 312938 345866 313174
rect 346102 312938 346134 313174
rect 345514 312854 346134 312938
rect 345514 312618 345546 312854
rect 345782 312618 345866 312854
rect 346102 312618 346134 312854
rect 345514 279174 346134 312618
rect 345514 278938 345546 279174
rect 345782 278938 345866 279174
rect 346102 278938 346134 279174
rect 345514 278854 346134 278938
rect 345514 278618 345546 278854
rect 345782 278618 345866 278854
rect 346102 278618 346134 278854
rect 345514 245174 346134 278618
rect 345514 244938 345546 245174
rect 345782 244938 345866 245174
rect 346102 244938 346134 245174
rect 345514 244854 346134 244938
rect 345514 244618 345546 244854
rect 345782 244618 345866 244854
rect 346102 244618 346134 244854
rect 345514 225660 346134 244618
rect 349234 706758 349854 711590
rect 349234 706522 349266 706758
rect 349502 706522 349586 706758
rect 349822 706522 349854 706758
rect 349234 706438 349854 706522
rect 349234 706202 349266 706438
rect 349502 706202 349586 706438
rect 349822 706202 349854 706438
rect 349234 690894 349854 706202
rect 349234 690658 349266 690894
rect 349502 690658 349586 690894
rect 349822 690658 349854 690894
rect 349234 690574 349854 690658
rect 349234 690338 349266 690574
rect 349502 690338 349586 690574
rect 349822 690338 349854 690574
rect 349234 656894 349854 690338
rect 349234 656658 349266 656894
rect 349502 656658 349586 656894
rect 349822 656658 349854 656894
rect 349234 656574 349854 656658
rect 349234 656338 349266 656574
rect 349502 656338 349586 656574
rect 349822 656338 349854 656574
rect 349234 622894 349854 656338
rect 349234 622658 349266 622894
rect 349502 622658 349586 622894
rect 349822 622658 349854 622894
rect 349234 622574 349854 622658
rect 349234 622338 349266 622574
rect 349502 622338 349586 622574
rect 349822 622338 349854 622574
rect 349234 588894 349854 622338
rect 349234 588658 349266 588894
rect 349502 588658 349586 588894
rect 349822 588658 349854 588894
rect 349234 588574 349854 588658
rect 349234 588338 349266 588574
rect 349502 588338 349586 588574
rect 349822 588338 349854 588574
rect 349234 554894 349854 588338
rect 349234 554658 349266 554894
rect 349502 554658 349586 554894
rect 349822 554658 349854 554894
rect 349234 554574 349854 554658
rect 349234 554338 349266 554574
rect 349502 554338 349586 554574
rect 349822 554338 349854 554574
rect 349234 520894 349854 554338
rect 349234 520658 349266 520894
rect 349502 520658 349586 520894
rect 349822 520658 349854 520894
rect 349234 520574 349854 520658
rect 349234 520338 349266 520574
rect 349502 520338 349586 520574
rect 349822 520338 349854 520574
rect 349234 486894 349854 520338
rect 349234 486658 349266 486894
rect 349502 486658 349586 486894
rect 349822 486658 349854 486894
rect 349234 486574 349854 486658
rect 349234 486338 349266 486574
rect 349502 486338 349586 486574
rect 349822 486338 349854 486574
rect 349234 452894 349854 486338
rect 349234 452658 349266 452894
rect 349502 452658 349586 452894
rect 349822 452658 349854 452894
rect 349234 452574 349854 452658
rect 349234 452338 349266 452574
rect 349502 452338 349586 452574
rect 349822 452338 349854 452574
rect 349234 418894 349854 452338
rect 349234 418658 349266 418894
rect 349502 418658 349586 418894
rect 349822 418658 349854 418894
rect 349234 418574 349854 418658
rect 349234 418338 349266 418574
rect 349502 418338 349586 418574
rect 349822 418338 349854 418574
rect 349234 384894 349854 418338
rect 349234 384658 349266 384894
rect 349502 384658 349586 384894
rect 349822 384658 349854 384894
rect 349234 384574 349854 384658
rect 349234 384338 349266 384574
rect 349502 384338 349586 384574
rect 349822 384338 349854 384574
rect 349234 350894 349854 384338
rect 349234 350658 349266 350894
rect 349502 350658 349586 350894
rect 349822 350658 349854 350894
rect 349234 350574 349854 350658
rect 349234 350338 349266 350574
rect 349502 350338 349586 350574
rect 349822 350338 349854 350574
rect 349234 316894 349854 350338
rect 349234 316658 349266 316894
rect 349502 316658 349586 316894
rect 349822 316658 349854 316894
rect 349234 316574 349854 316658
rect 349234 316338 349266 316574
rect 349502 316338 349586 316574
rect 349822 316338 349854 316574
rect 349234 282894 349854 316338
rect 349234 282658 349266 282894
rect 349502 282658 349586 282894
rect 349822 282658 349854 282894
rect 349234 282574 349854 282658
rect 349234 282338 349266 282574
rect 349502 282338 349586 282574
rect 349822 282338 349854 282574
rect 349234 248894 349854 282338
rect 349234 248658 349266 248894
rect 349502 248658 349586 248894
rect 349822 248658 349854 248894
rect 349234 248574 349854 248658
rect 349234 248338 349266 248574
rect 349502 248338 349586 248574
rect 349822 248338 349854 248574
rect 349234 225660 349854 248338
rect 352954 707718 353574 711590
rect 352954 707482 352986 707718
rect 353222 707482 353306 707718
rect 353542 707482 353574 707718
rect 352954 707398 353574 707482
rect 352954 707162 352986 707398
rect 353222 707162 353306 707398
rect 353542 707162 353574 707398
rect 352954 694614 353574 707162
rect 352954 694378 352986 694614
rect 353222 694378 353306 694614
rect 353542 694378 353574 694614
rect 352954 694294 353574 694378
rect 352954 694058 352986 694294
rect 353222 694058 353306 694294
rect 353542 694058 353574 694294
rect 352954 660614 353574 694058
rect 352954 660378 352986 660614
rect 353222 660378 353306 660614
rect 353542 660378 353574 660614
rect 352954 660294 353574 660378
rect 352954 660058 352986 660294
rect 353222 660058 353306 660294
rect 353542 660058 353574 660294
rect 352954 626614 353574 660058
rect 352954 626378 352986 626614
rect 353222 626378 353306 626614
rect 353542 626378 353574 626614
rect 352954 626294 353574 626378
rect 352954 626058 352986 626294
rect 353222 626058 353306 626294
rect 353542 626058 353574 626294
rect 352954 592614 353574 626058
rect 352954 592378 352986 592614
rect 353222 592378 353306 592614
rect 353542 592378 353574 592614
rect 352954 592294 353574 592378
rect 352954 592058 352986 592294
rect 353222 592058 353306 592294
rect 353542 592058 353574 592294
rect 352954 558614 353574 592058
rect 352954 558378 352986 558614
rect 353222 558378 353306 558614
rect 353542 558378 353574 558614
rect 352954 558294 353574 558378
rect 352954 558058 352986 558294
rect 353222 558058 353306 558294
rect 353542 558058 353574 558294
rect 352954 524614 353574 558058
rect 352954 524378 352986 524614
rect 353222 524378 353306 524614
rect 353542 524378 353574 524614
rect 352954 524294 353574 524378
rect 352954 524058 352986 524294
rect 353222 524058 353306 524294
rect 353542 524058 353574 524294
rect 352954 490614 353574 524058
rect 352954 490378 352986 490614
rect 353222 490378 353306 490614
rect 353542 490378 353574 490614
rect 352954 490294 353574 490378
rect 352954 490058 352986 490294
rect 353222 490058 353306 490294
rect 353542 490058 353574 490294
rect 352954 456614 353574 490058
rect 352954 456378 352986 456614
rect 353222 456378 353306 456614
rect 353542 456378 353574 456614
rect 352954 456294 353574 456378
rect 352954 456058 352986 456294
rect 353222 456058 353306 456294
rect 353542 456058 353574 456294
rect 352954 422614 353574 456058
rect 352954 422378 352986 422614
rect 353222 422378 353306 422614
rect 353542 422378 353574 422614
rect 352954 422294 353574 422378
rect 352954 422058 352986 422294
rect 353222 422058 353306 422294
rect 353542 422058 353574 422294
rect 352954 388614 353574 422058
rect 352954 388378 352986 388614
rect 353222 388378 353306 388614
rect 353542 388378 353574 388614
rect 352954 388294 353574 388378
rect 352954 388058 352986 388294
rect 353222 388058 353306 388294
rect 353542 388058 353574 388294
rect 352954 354614 353574 388058
rect 352954 354378 352986 354614
rect 353222 354378 353306 354614
rect 353542 354378 353574 354614
rect 352954 354294 353574 354378
rect 352954 354058 352986 354294
rect 353222 354058 353306 354294
rect 353542 354058 353574 354294
rect 352954 320614 353574 354058
rect 352954 320378 352986 320614
rect 353222 320378 353306 320614
rect 353542 320378 353574 320614
rect 352954 320294 353574 320378
rect 352954 320058 352986 320294
rect 353222 320058 353306 320294
rect 353542 320058 353574 320294
rect 352954 286614 353574 320058
rect 352954 286378 352986 286614
rect 353222 286378 353306 286614
rect 353542 286378 353574 286614
rect 352954 286294 353574 286378
rect 352954 286058 352986 286294
rect 353222 286058 353306 286294
rect 353542 286058 353574 286294
rect 352954 252614 353574 286058
rect 352954 252378 352986 252614
rect 353222 252378 353306 252614
rect 353542 252378 353574 252614
rect 352954 252294 353574 252378
rect 352954 252058 352986 252294
rect 353222 252058 353306 252294
rect 353542 252058 353574 252294
rect 352954 225660 353574 252058
rect 356674 708678 357294 711590
rect 356674 708442 356706 708678
rect 356942 708442 357026 708678
rect 357262 708442 357294 708678
rect 356674 708358 357294 708442
rect 356674 708122 356706 708358
rect 356942 708122 357026 708358
rect 357262 708122 357294 708358
rect 356674 698334 357294 708122
rect 356674 698098 356706 698334
rect 356942 698098 357026 698334
rect 357262 698098 357294 698334
rect 356674 698014 357294 698098
rect 356674 697778 356706 698014
rect 356942 697778 357026 698014
rect 357262 697778 357294 698014
rect 356674 664334 357294 697778
rect 356674 664098 356706 664334
rect 356942 664098 357026 664334
rect 357262 664098 357294 664334
rect 356674 664014 357294 664098
rect 356674 663778 356706 664014
rect 356942 663778 357026 664014
rect 357262 663778 357294 664014
rect 356674 630334 357294 663778
rect 356674 630098 356706 630334
rect 356942 630098 357026 630334
rect 357262 630098 357294 630334
rect 356674 630014 357294 630098
rect 356674 629778 356706 630014
rect 356942 629778 357026 630014
rect 357262 629778 357294 630014
rect 356674 596334 357294 629778
rect 356674 596098 356706 596334
rect 356942 596098 357026 596334
rect 357262 596098 357294 596334
rect 356674 596014 357294 596098
rect 356674 595778 356706 596014
rect 356942 595778 357026 596014
rect 357262 595778 357294 596014
rect 356674 562334 357294 595778
rect 356674 562098 356706 562334
rect 356942 562098 357026 562334
rect 357262 562098 357294 562334
rect 356674 562014 357294 562098
rect 356674 561778 356706 562014
rect 356942 561778 357026 562014
rect 357262 561778 357294 562014
rect 356674 528334 357294 561778
rect 356674 528098 356706 528334
rect 356942 528098 357026 528334
rect 357262 528098 357294 528334
rect 356674 528014 357294 528098
rect 356674 527778 356706 528014
rect 356942 527778 357026 528014
rect 357262 527778 357294 528014
rect 356674 494334 357294 527778
rect 356674 494098 356706 494334
rect 356942 494098 357026 494334
rect 357262 494098 357294 494334
rect 356674 494014 357294 494098
rect 356674 493778 356706 494014
rect 356942 493778 357026 494014
rect 357262 493778 357294 494014
rect 356674 460334 357294 493778
rect 356674 460098 356706 460334
rect 356942 460098 357026 460334
rect 357262 460098 357294 460334
rect 356674 460014 357294 460098
rect 356674 459778 356706 460014
rect 356942 459778 357026 460014
rect 357262 459778 357294 460014
rect 356674 426334 357294 459778
rect 356674 426098 356706 426334
rect 356942 426098 357026 426334
rect 357262 426098 357294 426334
rect 356674 426014 357294 426098
rect 356674 425778 356706 426014
rect 356942 425778 357026 426014
rect 357262 425778 357294 426014
rect 356674 392334 357294 425778
rect 356674 392098 356706 392334
rect 356942 392098 357026 392334
rect 357262 392098 357294 392334
rect 356674 392014 357294 392098
rect 356674 391778 356706 392014
rect 356942 391778 357026 392014
rect 357262 391778 357294 392014
rect 356674 358334 357294 391778
rect 356674 358098 356706 358334
rect 356942 358098 357026 358334
rect 357262 358098 357294 358334
rect 356674 358014 357294 358098
rect 356674 357778 356706 358014
rect 356942 357778 357026 358014
rect 357262 357778 357294 358014
rect 356674 324334 357294 357778
rect 356674 324098 356706 324334
rect 356942 324098 357026 324334
rect 357262 324098 357294 324334
rect 356674 324014 357294 324098
rect 356674 323778 356706 324014
rect 356942 323778 357026 324014
rect 357262 323778 357294 324014
rect 356674 290334 357294 323778
rect 356674 290098 356706 290334
rect 356942 290098 357026 290334
rect 357262 290098 357294 290334
rect 356674 290014 357294 290098
rect 356674 289778 356706 290014
rect 356942 289778 357026 290014
rect 357262 289778 357294 290014
rect 356674 256334 357294 289778
rect 356674 256098 356706 256334
rect 356942 256098 357026 256334
rect 357262 256098 357294 256334
rect 356674 256014 357294 256098
rect 356674 255778 356706 256014
rect 356942 255778 357026 256014
rect 357262 255778 357294 256014
rect 356674 225660 357294 255778
rect 360394 709638 361014 711590
rect 360394 709402 360426 709638
rect 360662 709402 360746 709638
rect 360982 709402 361014 709638
rect 360394 709318 361014 709402
rect 360394 709082 360426 709318
rect 360662 709082 360746 709318
rect 360982 709082 361014 709318
rect 360394 668054 361014 709082
rect 360394 667818 360426 668054
rect 360662 667818 360746 668054
rect 360982 667818 361014 668054
rect 360394 667734 361014 667818
rect 360394 667498 360426 667734
rect 360662 667498 360746 667734
rect 360982 667498 361014 667734
rect 360394 634054 361014 667498
rect 360394 633818 360426 634054
rect 360662 633818 360746 634054
rect 360982 633818 361014 634054
rect 360394 633734 361014 633818
rect 360394 633498 360426 633734
rect 360662 633498 360746 633734
rect 360982 633498 361014 633734
rect 360394 600054 361014 633498
rect 360394 599818 360426 600054
rect 360662 599818 360746 600054
rect 360982 599818 361014 600054
rect 360394 599734 361014 599818
rect 360394 599498 360426 599734
rect 360662 599498 360746 599734
rect 360982 599498 361014 599734
rect 360394 566054 361014 599498
rect 360394 565818 360426 566054
rect 360662 565818 360746 566054
rect 360982 565818 361014 566054
rect 360394 565734 361014 565818
rect 360394 565498 360426 565734
rect 360662 565498 360746 565734
rect 360982 565498 361014 565734
rect 360394 532054 361014 565498
rect 360394 531818 360426 532054
rect 360662 531818 360746 532054
rect 360982 531818 361014 532054
rect 360394 531734 361014 531818
rect 360394 531498 360426 531734
rect 360662 531498 360746 531734
rect 360982 531498 361014 531734
rect 360394 498054 361014 531498
rect 360394 497818 360426 498054
rect 360662 497818 360746 498054
rect 360982 497818 361014 498054
rect 360394 497734 361014 497818
rect 360394 497498 360426 497734
rect 360662 497498 360746 497734
rect 360982 497498 361014 497734
rect 360394 464054 361014 497498
rect 360394 463818 360426 464054
rect 360662 463818 360746 464054
rect 360982 463818 361014 464054
rect 360394 463734 361014 463818
rect 360394 463498 360426 463734
rect 360662 463498 360746 463734
rect 360982 463498 361014 463734
rect 360394 430054 361014 463498
rect 360394 429818 360426 430054
rect 360662 429818 360746 430054
rect 360982 429818 361014 430054
rect 360394 429734 361014 429818
rect 360394 429498 360426 429734
rect 360662 429498 360746 429734
rect 360982 429498 361014 429734
rect 360394 396054 361014 429498
rect 360394 395818 360426 396054
rect 360662 395818 360746 396054
rect 360982 395818 361014 396054
rect 360394 395734 361014 395818
rect 360394 395498 360426 395734
rect 360662 395498 360746 395734
rect 360982 395498 361014 395734
rect 360394 362054 361014 395498
rect 360394 361818 360426 362054
rect 360662 361818 360746 362054
rect 360982 361818 361014 362054
rect 360394 361734 361014 361818
rect 360394 361498 360426 361734
rect 360662 361498 360746 361734
rect 360982 361498 361014 361734
rect 360394 328054 361014 361498
rect 360394 327818 360426 328054
rect 360662 327818 360746 328054
rect 360982 327818 361014 328054
rect 360394 327734 361014 327818
rect 360394 327498 360426 327734
rect 360662 327498 360746 327734
rect 360982 327498 361014 327734
rect 360394 294054 361014 327498
rect 360394 293818 360426 294054
rect 360662 293818 360746 294054
rect 360982 293818 361014 294054
rect 360394 293734 361014 293818
rect 360394 293498 360426 293734
rect 360662 293498 360746 293734
rect 360982 293498 361014 293734
rect 360394 260054 361014 293498
rect 360394 259818 360426 260054
rect 360662 259818 360746 260054
rect 360982 259818 361014 260054
rect 360394 259734 361014 259818
rect 360394 259498 360426 259734
rect 360662 259498 360746 259734
rect 360982 259498 361014 259734
rect 360394 225991 361014 259498
rect 360394 225755 360426 225991
rect 360662 225755 360746 225991
rect 360982 225755 361014 225991
rect 360394 225660 361014 225755
rect 364114 710598 364734 711590
rect 364114 710362 364146 710598
rect 364382 710362 364466 710598
rect 364702 710362 364734 710598
rect 364114 710278 364734 710362
rect 364114 710042 364146 710278
rect 364382 710042 364466 710278
rect 364702 710042 364734 710278
rect 364114 671774 364734 710042
rect 364114 671538 364146 671774
rect 364382 671538 364466 671774
rect 364702 671538 364734 671774
rect 364114 671454 364734 671538
rect 364114 671218 364146 671454
rect 364382 671218 364466 671454
rect 364702 671218 364734 671454
rect 364114 637774 364734 671218
rect 364114 637538 364146 637774
rect 364382 637538 364466 637774
rect 364702 637538 364734 637774
rect 364114 637454 364734 637538
rect 364114 637218 364146 637454
rect 364382 637218 364466 637454
rect 364702 637218 364734 637454
rect 364114 603774 364734 637218
rect 364114 603538 364146 603774
rect 364382 603538 364466 603774
rect 364702 603538 364734 603774
rect 364114 603454 364734 603538
rect 364114 603218 364146 603454
rect 364382 603218 364466 603454
rect 364702 603218 364734 603454
rect 364114 569774 364734 603218
rect 364114 569538 364146 569774
rect 364382 569538 364466 569774
rect 364702 569538 364734 569774
rect 364114 569454 364734 569538
rect 364114 569218 364146 569454
rect 364382 569218 364466 569454
rect 364702 569218 364734 569454
rect 364114 535774 364734 569218
rect 364114 535538 364146 535774
rect 364382 535538 364466 535774
rect 364702 535538 364734 535774
rect 364114 535454 364734 535538
rect 364114 535218 364146 535454
rect 364382 535218 364466 535454
rect 364702 535218 364734 535454
rect 364114 501774 364734 535218
rect 364114 501538 364146 501774
rect 364382 501538 364466 501774
rect 364702 501538 364734 501774
rect 364114 501454 364734 501538
rect 364114 501218 364146 501454
rect 364382 501218 364466 501454
rect 364702 501218 364734 501454
rect 364114 467774 364734 501218
rect 364114 467538 364146 467774
rect 364382 467538 364466 467774
rect 364702 467538 364734 467774
rect 364114 467454 364734 467538
rect 364114 467218 364146 467454
rect 364382 467218 364466 467454
rect 364702 467218 364734 467454
rect 364114 433774 364734 467218
rect 364114 433538 364146 433774
rect 364382 433538 364466 433774
rect 364702 433538 364734 433774
rect 364114 433454 364734 433538
rect 364114 433218 364146 433454
rect 364382 433218 364466 433454
rect 364702 433218 364734 433454
rect 364114 399774 364734 433218
rect 364114 399538 364146 399774
rect 364382 399538 364466 399774
rect 364702 399538 364734 399774
rect 364114 399454 364734 399538
rect 364114 399218 364146 399454
rect 364382 399218 364466 399454
rect 364702 399218 364734 399454
rect 364114 365774 364734 399218
rect 364114 365538 364146 365774
rect 364382 365538 364466 365774
rect 364702 365538 364734 365774
rect 364114 365454 364734 365538
rect 364114 365218 364146 365454
rect 364382 365218 364466 365454
rect 364702 365218 364734 365454
rect 364114 331774 364734 365218
rect 364114 331538 364146 331774
rect 364382 331538 364466 331774
rect 364702 331538 364734 331774
rect 364114 331454 364734 331538
rect 364114 331218 364146 331454
rect 364382 331218 364466 331454
rect 364702 331218 364734 331454
rect 364114 297774 364734 331218
rect 364114 297538 364146 297774
rect 364382 297538 364466 297774
rect 364702 297538 364734 297774
rect 364114 297454 364734 297538
rect 364114 297218 364146 297454
rect 364382 297218 364466 297454
rect 364702 297218 364734 297454
rect 364114 263774 364734 297218
rect 364114 263538 364146 263774
rect 364382 263538 364466 263774
rect 364702 263538 364734 263774
rect 364114 263454 364734 263538
rect 364114 263218 364146 263454
rect 364382 263218 364466 263454
rect 364702 263218 364734 263454
rect 364114 229774 364734 263218
rect 364114 229538 364146 229774
rect 364382 229538 364466 229774
rect 364702 229538 364734 229774
rect 364114 229454 364734 229538
rect 364114 229218 364146 229454
rect 364382 229218 364466 229454
rect 364702 229218 364734 229454
rect 364114 225660 364734 229218
rect 367834 711558 368454 711590
rect 367834 711322 367866 711558
rect 368102 711322 368186 711558
rect 368422 711322 368454 711558
rect 367834 711238 368454 711322
rect 367834 711002 367866 711238
rect 368102 711002 368186 711238
rect 368422 711002 368454 711238
rect 367834 675494 368454 711002
rect 367834 675258 367866 675494
rect 368102 675258 368186 675494
rect 368422 675258 368454 675494
rect 367834 675174 368454 675258
rect 367834 674938 367866 675174
rect 368102 674938 368186 675174
rect 368422 674938 368454 675174
rect 367834 641494 368454 674938
rect 367834 641258 367866 641494
rect 368102 641258 368186 641494
rect 368422 641258 368454 641494
rect 367834 641174 368454 641258
rect 367834 640938 367866 641174
rect 368102 640938 368186 641174
rect 368422 640938 368454 641174
rect 367834 607494 368454 640938
rect 367834 607258 367866 607494
rect 368102 607258 368186 607494
rect 368422 607258 368454 607494
rect 367834 607174 368454 607258
rect 367834 606938 367866 607174
rect 368102 606938 368186 607174
rect 368422 606938 368454 607174
rect 367834 573494 368454 606938
rect 367834 573258 367866 573494
rect 368102 573258 368186 573494
rect 368422 573258 368454 573494
rect 367834 573174 368454 573258
rect 367834 572938 367866 573174
rect 368102 572938 368186 573174
rect 368422 572938 368454 573174
rect 367834 539494 368454 572938
rect 367834 539258 367866 539494
rect 368102 539258 368186 539494
rect 368422 539258 368454 539494
rect 367834 539174 368454 539258
rect 367834 538938 367866 539174
rect 368102 538938 368186 539174
rect 368422 538938 368454 539174
rect 367834 505494 368454 538938
rect 367834 505258 367866 505494
rect 368102 505258 368186 505494
rect 368422 505258 368454 505494
rect 367834 505174 368454 505258
rect 367834 504938 367866 505174
rect 368102 504938 368186 505174
rect 368422 504938 368454 505174
rect 367834 471494 368454 504938
rect 367834 471258 367866 471494
rect 368102 471258 368186 471494
rect 368422 471258 368454 471494
rect 367834 471174 368454 471258
rect 367834 470938 367866 471174
rect 368102 470938 368186 471174
rect 368422 470938 368454 471174
rect 367834 437494 368454 470938
rect 367834 437258 367866 437494
rect 368102 437258 368186 437494
rect 368422 437258 368454 437494
rect 367834 437174 368454 437258
rect 367834 436938 367866 437174
rect 368102 436938 368186 437174
rect 368422 436938 368454 437174
rect 367834 403494 368454 436938
rect 367834 403258 367866 403494
rect 368102 403258 368186 403494
rect 368422 403258 368454 403494
rect 367834 403174 368454 403258
rect 367834 402938 367866 403174
rect 368102 402938 368186 403174
rect 368422 402938 368454 403174
rect 367834 369494 368454 402938
rect 367834 369258 367866 369494
rect 368102 369258 368186 369494
rect 368422 369258 368454 369494
rect 367834 369174 368454 369258
rect 367834 368938 367866 369174
rect 368102 368938 368186 369174
rect 368422 368938 368454 369174
rect 367834 335494 368454 368938
rect 367834 335258 367866 335494
rect 368102 335258 368186 335494
rect 368422 335258 368454 335494
rect 367834 335174 368454 335258
rect 367834 334938 367866 335174
rect 368102 334938 368186 335174
rect 368422 334938 368454 335174
rect 367834 301494 368454 334938
rect 367834 301258 367866 301494
rect 368102 301258 368186 301494
rect 368422 301258 368454 301494
rect 367834 301174 368454 301258
rect 367834 300938 367866 301174
rect 368102 300938 368186 301174
rect 368422 300938 368454 301174
rect 367834 267494 368454 300938
rect 367834 267258 367866 267494
rect 368102 267258 368186 267494
rect 368422 267258 368454 267494
rect 367834 267174 368454 267258
rect 367834 266938 367866 267174
rect 368102 266938 368186 267174
rect 368422 266938 368454 267174
rect 367834 233494 368454 266938
rect 367834 233258 367866 233494
rect 368102 233258 368186 233494
rect 368422 233258 368454 233494
rect 367834 233174 368454 233258
rect 367834 232938 367866 233174
rect 368102 232938 368186 233174
rect 368422 232938 368454 233174
rect 367834 225660 368454 232938
rect 375794 704838 376414 711590
rect 375794 704602 375826 704838
rect 376062 704602 376146 704838
rect 376382 704602 376414 704838
rect 375794 704518 376414 704602
rect 375794 704282 375826 704518
rect 376062 704282 376146 704518
rect 376382 704282 376414 704518
rect 375794 683454 376414 704282
rect 375794 683218 375826 683454
rect 376062 683218 376146 683454
rect 376382 683218 376414 683454
rect 375794 683134 376414 683218
rect 375794 682898 375826 683134
rect 376062 682898 376146 683134
rect 376382 682898 376414 683134
rect 375794 649454 376414 682898
rect 375794 649218 375826 649454
rect 376062 649218 376146 649454
rect 376382 649218 376414 649454
rect 375794 649134 376414 649218
rect 375794 648898 375826 649134
rect 376062 648898 376146 649134
rect 376382 648898 376414 649134
rect 375794 615454 376414 648898
rect 375794 615218 375826 615454
rect 376062 615218 376146 615454
rect 376382 615218 376414 615454
rect 375794 615134 376414 615218
rect 375794 614898 375826 615134
rect 376062 614898 376146 615134
rect 376382 614898 376414 615134
rect 375794 581454 376414 614898
rect 375794 581218 375826 581454
rect 376062 581218 376146 581454
rect 376382 581218 376414 581454
rect 375794 581134 376414 581218
rect 375794 580898 375826 581134
rect 376062 580898 376146 581134
rect 376382 580898 376414 581134
rect 375794 547454 376414 580898
rect 375794 547218 375826 547454
rect 376062 547218 376146 547454
rect 376382 547218 376414 547454
rect 375794 547134 376414 547218
rect 375794 546898 375826 547134
rect 376062 546898 376146 547134
rect 376382 546898 376414 547134
rect 375794 513454 376414 546898
rect 375794 513218 375826 513454
rect 376062 513218 376146 513454
rect 376382 513218 376414 513454
rect 375794 513134 376414 513218
rect 375794 512898 375826 513134
rect 376062 512898 376146 513134
rect 376382 512898 376414 513134
rect 375794 479454 376414 512898
rect 375794 479218 375826 479454
rect 376062 479218 376146 479454
rect 376382 479218 376414 479454
rect 375794 479134 376414 479218
rect 375794 478898 375826 479134
rect 376062 478898 376146 479134
rect 376382 478898 376414 479134
rect 375794 445454 376414 478898
rect 375794 445218 375826 445454
rect 376062 445218 376146 445454
rect 376382 445218 376414 445454
rect 375794 445134 376414 445218
rect 375794 444898 375826 445134
rect 376062 444898 376146 445134
rect 376382 444898 376414 445134
rect 375794 411454 376414 444898
rect 375794 411218 375826 411454
rect 376062 411218 376146 411454
rect 376382 411218 376414 411454
rect 375794 411134 376414 411218
rect 375794 410898 375826 411134
rect 376062 410898 376146 411134
rect 376382 410898 376414 411134
rect 375794 377454 376414 410898
rect 375794 377218 375826 377454
rect 376062 377218 376146 377454
rect 376382 377218 376414 377454
rect 375794 377134 376414 377218
rect 375794 376898 375826 377134
rect 376062 376898 376146 377134
rect 376382 376898 376414 377134
rect 375794 343454 376414 376898
rect 375794 343218 375826 343454
rect 376062 343218 376146 343454
rect 376382 343218 376414 343454
rect 375794 343134 376414 343218
rect 375794 342898 375826 343134
rect 376062 342898 376146 343134
rect 376382 342898 376414 343134
rect 375794 309454 376414 342898
rect 375794 309218 375826 309454
rect 376062 309218 376146 309454
rect 376382 309218 376414 309454
rect 375794 309134 376414 309218
rect 375794 308898 375826 309134
rect 376062 308898 376146 309134
rect 376382 308898 376414 309134
rect 375794 275454 376414 308898
rect 375794 275218 375826 275454
rect 376062 275218 376146 275454
rect 376382 275218 376414 275454
rect 375794 275134 376414 275218
rect 375794 274898 375826 275134
rect 376062 274898 376146 275134
rect 376382 274898 376414 275134
rect 375794 241454 376414 274898
rect 375794 241218 375826 241454
rect 376062 241218 376146 241454
rect 376382 241218 376414 241454
rect 375794 241134 376414 241218
rect 375794 240898 375826 241134
rect 376062 240898 376146 241134
rect 376382 240898 376414 241134
rect 375794 225660 376414 240898
rect 379514 705798 380134 711590
rect 379514 705562 379546 705798
rect 379782 705562 379866 705798
rect 380102 705562 380134 705798
rect 379514 705478 380134 705562
rect 379514 705242 379546 705478
rect 379782 705242 379866 705478
rect 380102 705242 380134 705478
rect 379514 687174 380134 705242
rect 379514 686938 379546 687174
rect 379782 686938 379866 687174
rect 380102 686938 380134 687174
rect 379514 686854 380134 686938
rect 379514 686618 379546 686854
rect 379782 686618 379866 686854
rect 380102 686618 380134 686854
rect 379514 653174 380134 686618
rect 379514 652938 379546 653174
rect 379782 652938 379866 653174
rect 380102 652938 380134 653174
rect 379514 652854 380134 652938
rect 379514 652618 379546 652854
rect 379782 652618 379866 652854
rect 380102 652618 380134 652854
rect 379514 619174 380134 652618
rect 379514 618938 379546 619174
rect 379782 618938 379866 619174
rect 380102 618938 380134 619174
rect 379514 618854 380134 618938
rect 379514 618618 379546 618854
rect 379782 618618 379866 618854
rect 380102 618618 380134 618854
rect 379514 585174 380134 618618
rect 379514 584938 379546 585174
rect 379782 584938 379866 585174
rect 380102 584938 380134 585174
rect 379514 584854 380134 584938
rect 379514 584618 379546 584854
rect 379782 584618 379866 584854
rect 380102 584618 380134 584854
rect 379514 551174 380134 584618
rect 379514 550938 379546 551174
rect 379782 550938 379866 551174
rect 380102 550938 380134 551174
rect 379514 550854 380134 550938
rect 379514 550618 379546 550854
rect 379782 550618 379866 550854
rect 380102 550618 380134 550854
rect 379514 517174 380134 550618
rect 379514 516938 379546 517174
rect 379782 516938 379866 517174
rect 380102 516938 380134 517174
rect 379514 516854 380134 516938
rect 379514 516618 379546 516854
rect 379782 516618 379866 516854
rect 380102 516618 380134 516854
rect 379514 483174 380134 516618
rect 379514 482938 379546 483174
rect 379782 482938 379866 483174
rect 380102 482938 380134 483174
rect 379514 482854 380134 482938
rect 379514 482618 379546 482854
rect 379782 482618 379866 482854
rect 380102 482618 380134 482854
rect 379514 449174 380134 482618
rect 379514 448938 379546 449174
rect 379782 448938 379866 449174
rect 380102 448938 380134 449174
rect 379514 448854 380134 448938
rect 379514 448618 379546 448854
rect 379782 448618 379866 448854
rect 380102 448618 380134 448854
rect 379514 415174 380134 448618
rect 379514 414938 379546 415174
rect 379782 414938 379866 415174
rect 380102 414938 380134 415174
rect 379514 414854 380134 414938
rect 379514 414618 379546 414854
rect 379782 414618 379866 414854
rect 380102 414618 380134 414854
rect 379514 381174 380134 414618
rect 379514 380938 379546 381174
rect 379782 380938 379866 381174
rect 380102 380938 380134 381174
rect 379514 380854 380134 380938
rect 379514 380618 379546 380854
rect 379782 380618 379866 380854
rect 380102 380618 380134 380854
rect 379514 347174 380134 380618
rect 379514 346938 379546 347174
rect 379782 346938 379866 347174
rect 380102 346938 380134 347174
rect 379514 346854 380134 346938
rect 379514 346618 379546 346854
rect 379782 346618 379866 346854
rect 380102 346618 380134 346854
rect 379514 313174 380134 346618
rect 379514 312938 379546 313174
rect 379782 312938 379866 313174
rect 380102 312938 380134 313174
rect 379514 312854 380134 312938
rect 379514 312618 379546 312854
rect 379782 312618 379866 312854
rect 380102 312618 380134 312854
rect 379514 279174 380134 312618
rect 379514 278938 379546 279174
rect 379782 278938 379866 279174
rect 380102 278938 380134 279174
rect 379514 278854 380134 278938
rect 379514 278618 379546 278854
rect 379782 278618 379866 278854
rect 380102 278618 380134 278854
rect 379514 245174 380134 278618
rect 379514 244938 379546 245174
rect 379782 244938 379866 245174
rect 380102 244938 380134 245174
rect 379514 244854 380134 244938
rect 379514 244618 379546 244854
rect 379782 244618 379866 244854
rect 380102 244618 380134 244854
rect 379514 225660 380134 244618
rect 383234 706758 383854 711590
rect 383234 706522 383266 706758
rect 383502 706522 383586 706758
rect 383822 706522 383854 706758
rect 383234 706438 383854 706522
rect 383234 706202 383266 706438
rect 383502 706202 383586 706438
rect 383822 706202 383854 706438
rect 383234 690894 383854 706202
rect 383234 690658 383266 690894
rect 383502 690658 383586 690894
rect 383822 690658 383854 690894
rect 383234 690574 383854 690658
rect 383234 690338 383266 690574
rect 383502 690338 383586 690574
rect 383822 690338 383854 690574
rect 383234 656894 383854 690338
rect 383234 656658 383266 656894
rect 383502 656658 383586 656894
rect 383822 656658 383854 656894
rect 383234 656574 383854 656658
rect 383234 656338 383266 656574
rect 383502 656338 383586 656574
rect 383822 656338 383854 656574
rect 383234 622894 383854 656338
rect 383234 622658 383266 622894
rect 383502 622658 383586 622894
rect 383822 622658 383854 622894
rect 383234 622574 383854 622658
rect 383234 622338 383266 622574
rect 383502 622338 383586 622574
rect 383822 622338 383854 622574
rect 383234 588894 383854 622338
rect 383234 588658 383266 588894
rect 383502 588658 383586 588894
rect 383822 588658 383854 588894
rect 383234 588574 383854 588658
rect 383234 588338 383266 588574
rect 383502 588338 383586 588574
rect 383822 588338 383854 588574
rect 383234 554894 383854 588338
rect 383234 554658 383266 554894
rect 383502 554658 383586 554894
rect 383822 554658 383854 554894
rect 383234 554574 383854 554658
rect 383234 554338 383266 554574
rect 383502 554338 383586 554574
rect 383822 554338 383854 554574
rect 383234 520894 383854 554338
rect 383234 520658 383266 520894
rect 383502 520658 383586 520894
rect 383822 520658 383854 520894
rect 383234 520574 383854 520658
rect 383234 520338 383266 520574
rect 383502 520338 383586 520574
rect 383822 520338 383854 520574
rect 383234 486894 383854 520338
rect 383234 486658 383266 486894
rect 383502 486658 383586 486894
rect 383822 486658 383854 486894
rect 383234 486574 383854 486658
rect 383234 486338 383266 486574
rect 383502 486338 383586 486574
rect 383822 486338 383854 486574
rect 383234 452894 383854 486338
rect 383234 452658 383266 452894
rect 383502 452658 383586 452894
rect 383822 452658 383854 452894
rect 383234 452574 383854 452658
rect 383234 452338 383266 452574
rect 383502 452338 383586 452574
rect 383822 452338 383854 452574
rect 383234 418894 383854 452338
rect 383234 418658 383266 418894
rect 383502 418658 383586 418894
rect 383822 418658 383854 418894
rect 383234 418574 383854 418658
rect 383234 418338 383266 418574
rect 383502 418338 383586 418574
rect 383822 418338 383854 418574
rect 383234 384894 383854 418338
rect 383234 384658 383266 384894
rect 383502 384658 383586 384894
rect 383822 384658 383854 384894
rect 383234 384574 383854 384658
rect 383234 384338 383266 384574
rect 383502 384338 383586 384574
rect 383822 384338 383854 384574
rect 383234 350894 383854 384338
rect 383234 350658 383266 350894
rect 383502 350658 383586 350894
rect 383822 350658 383854 350894
rect 383234 350574 383854 350658
rect 383234 350338 383266 350574
rect 383502 350338 383586 350574
rect 383822 350338 383854 350574
rect 383234 316894 383854 350338
rect 383234 316658 383266 316894
rect 383502 316658 383586 316894
rect 383822 316658 383854 316894
rect 383234 316574 383854 316658
rect 383234 316338 383266 316574
rect 383502 316338 383586 316574
rect 383822 316338 383854 316574
rect 383234 282894 383854 316338
rect 383234 282658 383266 282894
rect 383502 282658 383586 282894
rect 383822 282658 383854 282894
rect 383234 282574 383854 282658
rect 383234 282338 383266 282574
rect 383502 282338 383586 282574
rect 383822 282338 383854 282574
rect 383234 248894 383854 282338
rect 383234 248658 383266 248894
rect 383502 248658 383586 248894
rect 383822 248658 383854 248894
rect 383234 248574 383854 248658
rect 383234 248338 383266 248574
rect 383502 248338 383586 248574
rect 383822 248338 383854 248574
rect 383234 225660 383854 248338
rect 386954 707718 387574 711590
rect 386954 707482 386986 707718
rect 387222 707482 387306 707718
rect 387542 707482 387574 707718
rect 386954 707398 387574 707482
rect 386954 707162 386986 707398
rect 387222 707162 387306 707398
rect 387542 707162 387574 707398
rect 386954 694614 387574 707162
rect 386954 694378 386986 694614
rect 387222 694378 387306 694614
rect 387542 694378 387574 694614
rect 386954 694294 387574 694378
rect 386954 694058 386986 694294
rect 387222 694058 387306 694294
rect 387542 694058 387574 694294
rect 386954 660614 387574 694058
rect 386954 660378 386986 660614
rect 387222 660378 387306 660614
rect 387542 660378 387574 660614
rect 386954 660294 387574 660378
rect 386954 660058 386986 660294
rect 387222 660058 387306 660294
rect 387542 660058 387574 660294
rect 386954 626614 387574 660058
rect 386954 626378 386986 626614
rect 387222 626378 387306 626614
rect 387542 626378 387574 626614
rect 386954 626294 387574 626378
rect 386954 626058 386986 626294
rect 387222 626058 387306 626294
rect 387542 626058 387574 626294
rect 386954 592614 387574 626058
rect 386954 592378 386986 592614
rect 387222 592378 387306 592614
rect 387542 592378 387574 592614
rect 386954 592294 387574 592378
rect 386954 592058 386986 592294
rect 387222 592058 387306 592294
rect 387542 592058 387574 592294
rect 386954 558614 387574 592058
rect 386954 558378 386986 558614
rect 387222 558378 387306 558614
rect 387542 558378 387574 558614
rect 386954 558294 387574 558378
rect 386954 558058 386986 558294
rect 387222 558058 387306 558294
rect 387542 558058 387574 558294
rect 386954 524614 387574 558058
rect 386954 524378 386986 524614
rect 387222 524378 387306 524614
rect 387542 524378 387574 524614
rect 386954 524294 387574 524378
rect 386954 524058 386986 524294
rect 387222 524058 387306 524294
rect 387542 524058 387574 524294
rect 386954 490614 387574 524058
rect 386954 490378 386986 490614
rect 387222 490378 387306 490614
rect 387542 490378 387574 490614
rect 386954 490294 387574 490378
rect 386954 490058 386986 490294
rect 387222 490058 387306 490294
rect 387542 490058 387574 490294
rect 386954 456614 387574 490058
rect 386954 456378 386986 456614
rect 387222 456378 387306 456614
rect 387542 456378 387574 456614
rect 386954 456294 387574 456378
rect 386954 456058 386986 456294
rect 387222 456058 387306 456294
rect 387542 456058 387574 456294
rect 386954 422614 387574 456058
rect 386954 422378 386986 422614
rect 387222 422378 387306 422614
rect 387542 422378 387574 422614
rect 386954 422294 387574 422378
rect 386954 422058 386986 422294
rect 387222 422058 387306 422294
rect 387542 422058 387574 422294
rect 386954 388614 387574 422058
rect 386954 388378 386986 388614
rect 387222 388378 387306 388614
rect 387542 388378 387574 388614
rect 386954 388294 387574 388378
rect 386954 388058 386986 388294
rect 387222 388058 387306 388294
rect 387542 388058 387574 388294
rect 386954 354614 387574 388058
rect 386954 354378 386986 354614
rect 387222 354378 387306 354614
rect 387542 354378 387574 354614
rect 386954 354294 387574 354378
rect 386954 354058 386986 354294
rect 387222 354058 387306 354294
rect 387542 354058 387574 354294
rect 386954 320614 387574 354058
rect 386954 320378 386986 320614
rect 387222 320378 387306 320614
rect 387542 320378 387574 320614
rect 386954 320294 387574 320378
rect 386954 320058 386986 320294
rect 387222 320058 387306 320294
rect 387542 320058 387574 320294
rect 386954 286614 387574 320058
rect 386954 286378 386986 286614
rect 387222 286378 387306 286614
rect 387542 286378 387574 286614
rect 386954 286294 387574 286378
rect 386954 286058 386986 286294
rect 387222 286058 387306 286294
rect 387542 286058 387574 286294
rect 386954 252614 387574 286058
rect 386954 252378 386986 252614
rect 387222 252378 387306 252614
rect 387542 252378 387574 252614
rect 386954 252294 387574 252378
rect 386954 252058 386986 252294
rect 387222 252058 387306 252294
rect 387542 252058 387574 252294
rect 386954 225660 387574 252058
rect 390674 708678 391294 711590
rect 390674 708442 390706 708678
rect 390942 708442 391026 708678
rect 391262 708442 391294 708678
rect 390674 708358 391294 708442
rect 390674 708122 390706 708358
rect 390942 708122 391026 708358
rect 391262 708122 391294 708358
rect 390674 698334 391294 708122
rect 390674 698098 390706 698334
rect 390942 698098 391026 698334
rect 391262 698098 391294 698334
rect 390674 698014 391294 698098
rect 390674 697778 390706 698014
rect 390942 697778 391026 698014
rect 391262 697778 391294 698014
rect 390674 664334 391294 697778
rect 390674 664098 390706 664334
rect 390942 664098 391026 664334
rect 391262 664098 391294 664334
rect 390674 664014 391294 664098
rect 390674 663778 390706 664014
rect 390942 663778 391026 664014
rect 391262 663778 391294 664014
rect 390674 630334 391294 663778
rect 390674 630098 390706 630334
rect 390942 630098 391026 630334
rect 391262 630098 391294 630334
rect 390674 630014 391294 630098
rect 390674 629778 390706 630014
rect 390942 629778 391026 630014
rect 391262 629778 391294 630014
rect 390674 596334 391294 629778
rect 390674 596098 390706 596334
rect 390942 596098 391026 596334
rect 391262 596098 391294 596334
rect 390674 596014 391294 596098
rect 390674 595778 390706 596014
rect 390942 595778 391026 596014
rect 391262 595778 391294 596014
rect 390674 562334 391294 595778
rect 390674 562098 390706 562334
rect 390942 562098 391026 562334
rect 391262 562098 391294 562334
rect 390674 562014 391294 562098
rect 390674 561778 390706 562014
rect 390942 561778 391026 562014
rect 391262 561778 391294 562014
rect 390674 528334 391294 561778
rect 390674 528098 390706 528334
rect 390942 528098 391026 528334
rect 391262 528098 391294 528334
rect 390674 528014 391294 528098
rect 390674 527778 390706 528014
rect 390942 527778 391026 528014
rect 391262 527778 391294 528014
rect 390674 494334 391294 527778
rect 390674 494098 390706 494334
rect 390942 494098 391026 494334
rect 391262 494098 391294 494334
rect 390674 494014 391294 494098
rect 390674 493778 390706 494014
rect 390942 493778 391026 494014
rect 391262 493778 391294 494014
rect 390674 460334 391294 493778
rect 390674 460098 390706 460334
rect 390942 460098 391026 460334
rect 391262 460098 391294 460334
rect 390674 460014 391294 460098
rect 390674 459778 390706 460014
rect 390942 459778 391026 460014
rect 391262 459778 391294 460014
rect 390674 426334 391294 459778
rect 390674 426098 390706 426334
rect 390942 426098 391026 426334
rect 391262 426098 391294 426334
rect 390674 426014 391294 426098
rect 390674 425778 390706 426014
rect 390942 425778 391026 426014
rect 391262 425778 391294 426014
rect 390674 392334 391294 425778
rect 390674 392098 390706 392334
rect 390942 392098 391026 392334
rect 391262 392098 391294 392334
rect 390674 392014 391294 392098
rect 390674 391778 390706 392014
rect 390942 391778 391026 392014
rect 391262 391778 391294 392014
rect 390674 358334 391294 391778
rect 390674 358098 390706 358334
rect 390942 358098 391026 358334
rect 391262 358098 391294 358334
rect 390674 358014 391294 358098
rect 390674 357778 390706 358014
rect 390942 357778 391026 358014
rect 391262 357778 391294 358014
rect 390674 324334 391294 357778
rect 390674 324098 390706 324334
rect 390942 324098 391026 324334
rect 391262 324098 391294 324334
rect 390674 324014 391294 324098
rect 390674 323778 390706 324014
rect 390942 323778 391026 324014
rect 391262 323778 391294 324014
rect 390674 290334 391294 323778
rect 390674 290098 390706 290334
rect 390942 290098 391026 290334
rect 391262 290098 391294 290334
rect 390674 290014 391294 290098
rect 390674 289778 390706 290014
rect 390942 289778 391026 290014
rect 391262 289778 391294 290014
rect 390674 256334 391294 289778
rect 390674 256098 390706 256334
rect 390942 256098 391026 256334
rect 391262 256098 391294 256334
rect 390674 256014 391294 256098
rect 390674 255778 390706 256014
rect 390942 255778 391026 256014
rect 391262 255778 391294 256014
rect 390674 225660 391294 255778
rect 394394 709638 395014 711590
rect 394394 709402 394426 709638
rect 394662 709402 394746 709638
rect 394982 709402 395014 709638
rect 394394 709318 395014 709402
rect 394394 709082 394426 709318
rect 394662 709082 394746 709318
rect 394982 709082 395014 709318
rect 394394 668054 395014 709082
rect 394394 667818 394426 668054
rect 394662 667818 394746 668054
rect 394982 667818 395014 668054
rect 394394 667734 395014 667818
rect 394394 667498 394426 667734
rect 394662 667498 394746 667734
rect 394982 667498 395014 667734
rect 394394 634054 395014 667498
rect 394394 633818 394426 634054
rect 394662 633818 394746 634054
rect 394982 633818 395014 634054
rect 394394 633734 395014 633818
rect 394394 633498 394426 633734
rect 394662 633498 394746 633734
rect 394982 633498 395014 633734
rect 394394 600054 395014 633498
rect 394394 599818 394426 600054
rect 394662 599818 394746 600054
rect 394982 599818 395014 600054
rect 394394 599734 395014 599818
rect 394394 599498 394426 599734
rect 394662 599498 394746 599734
rect 394982 599498 395014 599734
rect 394394 566054 395014 599498
rect 394394 565818 394426 566054
rect 394662 565818 394746 566054
rect 394982 565818 395014 566054
rect 394394 565734 395014 565818
rect 394394 565498 394426 565734
rect 394662 565498 394746 565734
rect 394982 565498 395014 565734
rect 394394 532054 395014 565498
rect 394394 531818 394426 532054
rect 394662 531818 394746 532054
rect 394982 531818 395014 532054
rect 394394 531734 395014 531818
rect 394394 531498 394426 531734
rect 394662 531498 394746 531734
rect 394982 531498 395014 531734
rect 394394 498054 395014 531498
rect 394394 497818 394426 498054
rect 394662 497818 394746 498054
rect 394982 497818 395014 498054
rect 394394 497734 395014 497818
rect 394394 497498 394426 497734
rect 394662 497498 394746 497734
rect 394982 497498 395014 497734
rect 394394 464054 395014 497498
rect 394394 463818 394426 464054
rect 394662 463818 394746 464054
rect 394982 463818 395014 464054
rect 394394 463734 395014 463818
rect 394394 463498 394426 463734
rect 394662 463498 394746 463734
rect 394982 463498 395014 463734
rect 394394 430054 395014 463498
rect 394394 429818 394426 430054
rect 394662 429818 394746 430054
rect 394982 429818 395014 430054
rect 394394 429734 395014 429818
rect 394394 429498 394426 429734
rect 394662 429498 394746 429734
rect 394982 429498 395014 429734
rect 394394 396054 395014 429498
rect 394394 395818 394426 396054
rect 394662 395818 394746 396054
rect 394982 395818 395014 396054
rect 394394 395734 395014 395818
rect 394394 395498 394426 395734
rect 394662 395498 394746 395734
rect 394982 395498 395014 395734
rect 394394 362054 395014 395498
rect 394394 361818 394426 362054
rect 394662 361818 394746 362054
rect 394982 361818 395014 362054
rect 394394 361734 395014 361818
rect 394394 361498 394426 361734
rect 394662 361498 394746 361734
rect 394982 361498 395014 361734
rect 394394 328054 395014 361498
rect 394394 327818 394426 328054
rect 394662 327818 394746 328054
rect 394982 327818 395014 328054
rect 394394 327734 395014 327818
rect 394394 327498 394426 327734
rect 394662 327498 394746 327734
rect 394982 327498 395014 327734
rect 394394 294054 395014 327498
rect 394394 293818 394426 294054
rect 394662 293818 394746 294054
rect 394982 293818 395014 294054
rect 394394 293734 395014 293818
rect 394394 293498 394426 293734
rect 394662 293498 394746 293734
rect 394982 293498 395014 293734
rect 394394 260054 395014 293498
rect 394394 259818 394426 260054
rect 394662 259818 394746 260054
rect 394982 259818 395014 260054
rect 394394 259734 395014 259818
rect 394394 259498 394426 259734
rect 394662 259498 394746 259734
rect 394982 259498 395014 259734
rect 394394 225991 395014 259498
rect 394394 225755 394426 225991
rect 394662 225755 394746 225991
rect 394982 225755 395014 225991
rect 394394 225660 395014 225755
rect 398114 710598 398734 711590
rect 398114 710362 398146 710598
rect 398382 710362 398466 710598
rect 398702 710362 398734 710598
rect 398114 710278 398734 710362
rect 398114 710042 398146 710278
rect 398382 710042 398466 710278
rect 398702 710042 398734 710278
rect 398114 671774 398734 710042
rect 398114 671538 398146 671774
rect 398382 671538 398466 671774
rect 398702 671538 398734 671774
rect 398114 671454 398734 671538
rect 398114 671218 398146 671454
rect 398382 671218 398466 671454
rect 398702 671218 398734 671454
rect 398114 637774 398734 671218
rect 398114 637538 398146 637774
rect 398382 637538 398466 637774
rect 398702 637538 398734 637774
rect 398114 637454 398734 637538
rect 398114 637218 398146 637454
rect 398382 637218 398466 637454
rect 398702 637218 398734 637454
rect 398114 603774 398734 637218
rect 398114 603538 398146 603774
rect 398382 603538 398466 603774
rect 398702 603538 398734 603774
rect 398114 603454 398734 603538
rect 398114 603218 398146 603454
rect 398382 603218 398466 603454
rect 398702 603218 398734 603454
rect 398114 569774 398734 603218
rect 398114 569538 398146 569774
rect 398382 569538 398466 569774
rect 398702 569538 398734 569774
rect 398114 569454 398734 569538
rect 398114 569218 398146 569454
rect 398382 569218 398466 569454
rect 398702 569218 398734 569454
rect 398114 535774 398734 569218
rect 398114 535538 398146 535774
rect 398382 535538 398466 535774
rect 398702 535538 398734 535774
rect 398114 535454 398734 535538
rect 398114 535218 398146 535454
rect 398382 535218 398466 535454
rect 398702 535218 398734 535454
rect 398114 501774 398734 535218
rect 398114 501538 398146 501774
rect 398382 501538 398466 501774
rect 398702 501538 398734 501774
rect 398114 501454 398734 501538
rect 398114 501218 398146 501454
rect 398382 501218 398466 501454
rect 398702 501218 398734 501454
rect 398114 467774 398734 501218
rect 398114 467538 398146 467774
rect 398382 467538 398466 467774
rect 398702 467538 398734 467774
rect 398114 467454 398734 467538
rect 398114 467218 398146 467454
rect 398382 467218 398466 467454
rect 398702 467218 398734 467454
rect 398114 433774 398734 467218
rect 398114 433538 398146 433774
rect 398382 433538 398466 433774
rect 398702 433538 398734 433774
rect 398114 433454 398734 433538
rect 398114 433218 398146 433454
rect 398382 433218 398466 433454
rect 398702 433218 398734 433454
rect 398114 399774 398734 433218
rect 398114 399538 398146 399774
rect 398382 399538 398466 399774
rect 398702 399538 398734 399774
rect 398114 399454 398734 399538
rect 398114 399218 398146 399454
rect 398382 399218 398466 399454
rect 398702 399218 398734 399454
rect 398114 365774 398734 399218
rect 398114 365538 398146 365774
rect 398382 365538 398466 365774
rect 398702 365538 398734 365774
rect 398114 365454 398734 365538
rect 398114 365218 398146 365454
rect 398382 365218 398466 365454
rect 398702 365218 398734 365454
rect 398114 331774 398734 365218
rect 398114 331538 398146 331774
rect 398382 331538 398466 331774
rect 398702 331538 398734 331774
rect 398114 331454 398734 331538
rect 398114 331218 398146 331454
rect 398382 331218 398466 331454
rect 398702 331218 398734 331454
rect 398114 297774 398734 331218
rect 398114 297538 398146 297774
rect 398382 297538 398466 297774
rect 398702 297538 398734 297774
rect 398114 297454 398734 297538
rect 398114 297218 398146 297454
rect 398382 297218 398466 297454
rect 398702 297218 398734 297454
rect 398114 263774 398734 297218
rect 398114 263538 398146 263774
rect 398382 263538 398466 263774
rect 398702 263538 398734 263774
rect 398114 263454 398734 263538
rect 398114 263218 398146 263454
rect 398382 263218 398466 263454
rect 398702 263218 398734 263454
rect 398114 229774 398734 263218
rect 398114 229538 398146 229774
rect 398382 229538 398466 229774
rect 398702 229538 398734 229774
rect 398114 229454 398734 229538
rect 398114 229218 398146 229454
rect 398382 229218 398466 229454
rect 398702 229218 398734 229454
rect 398114 225660 398734 229218
rect 401834 711558 402454 711590
rect 401834 711322 401866 711558
rect 402102 711322 402186 711558
rect 402422 711322 402454 711558
rect 401834 711238 402454 711322
rect 401834 711002 401866 711238
rect 402102 711002 402186 711238
rect 402422 711002 402454 711238
rect 401834 675494 402454 711002
rect 401834 675258 401866 675494
rect 402102 675258 402186 675494
rect 402422 675258 402454 675494
rect 401834 675174 402454 675258
rect 401834 674938 401866 675174
rect 402102 674938 402186 675174
rect 402422 674938 402454 675174
rect 401834 641494 402454 674938
rect 401834 641258 401866 641494
rect 402102 641258 402186 641494
rect 402422 641258 402454 641494
rect 401834 641174 402454 641258
rect 401834 640938 401866 641174
rect 402102 640938 402186 641174
rect 402422 640938 402454 641174
rect 401834 607494 402454 640938
rect 401834 607258 401866 607494
rect 402102 607258 402186 607494
rect 402422 607258 402454 607494
rect 401834 607174 402454 607258
rect 401834 606938 401866 607174
rect 402102 606938 402186 607174
rect 402422 606938 402454 607174
rect 401834 573494 402454 606938
rect 401834 573258 401866 573494
rect 402102 573258 402186 573494
rect 402422 573258 402454 573494
rect 401834 573174 402454 573258
rect 401834 572938 401866 573174
rect 402102 572938 402186 573174
rect 402422 572938 402454 573174
rect 401834 539494 402454 572938
rect 401834 539258 401866 539494
rect 402102 539258 402186 539494
rect 402422 539258 402454 539494
rect 401834 539174 402454 539258
rect 401834 538938 401866 539174
rect 402102 538938 402186 539174
rect 402422 538938 402454 539174
rect 401834 505494 402454 538938
rect 401834 505258 401866 505494
rect 402102 505258 402186 505494
rect 402422 505258 402454 505494
rect 401834 505174 402454 505258
rect 401834 504938 401866 505174
rect 402102 504938 402186 505174
rect 402422 504938 402454 505174
rect 401834 471494 402454 504938
rect 401834 471258 401866 471494
rect 402102 471258 402186 471494
rect 402422 471258 402454 471494
rect 401834 471174 402454 471258
rect 401834 470938 401866 471174
rect 402102 470938 402186 471174
rect 402422 470938 402454 471174
rect 401834 437494 402454 470938
rect 401834 437258 401866 437494
rect 402102 437258 402186 437494
rect 402422 437258 402454 437494
rect 401834 437174 402454 437258
rect 401834 436938 401866 437174
rect 402102 436938 402186 437174
rect 402422 436938 402454 437174
rect 401834 403494 402454 436938
rect 401834 403258 401866 403494
rect 402102 403258 402186 403494
rect 402422 403258 402454 403494
rect 401834 403174 402454 403258
rect 401834 402938 401866 403174
rect 402102 402938 402186 403174
rect 402422 402938 402454 403174
rect 401834 369494 402454 402938
rect 401834 369258 401866 369494
rect 402102 369258 402186 369494
rect 402422 369258 402454 369494
rect 401834 369174 402454 369258
rect 401834 368938 401866 369174
rect 402102 368938 402186 369174
rect 402422 368938 402454 369174
rect 401834 335494 402454 368938
rect 401834 335258 401866 335494
rect 402102 335258 402186 335494
rect 402422 335258 402454 335494
rect 401834 335174 402454 335258
rect 401834 334938 401866 335174
rect 402102 334938 402186 335174
rect 402422 334938 402454 335174
rect 401834 301494 402454 334938
rect 401834 301258 401866 301494
rect 402102 301258 402186 301494
rect 402422 301258 402454 301494
rect 401834 301174 402454 301258
rect 401834 300938 401866 301174
rect 402102 300938 402186 301174
rect 402422 300938 402454 301174
rect 401834 267494 402454 300938
rect 401834 267258 401866 267494
rect 402102 267258 402186 267494
rect 402422 267258 402454 267494
rect 401834 267174 402454 267258
rect 401834 266938 401866 267174
rect 402102 266938 402186 267174
rect 402422 266938 402454 267174
rect 401834 233494 402454 266938
rect 401834 233258 401866 233494
rect 402102 233258 402186 233494
rect 402422 233258 402454 233494
rect 401834 233174 402454 233258
rect 401834 232938 401866 233174
rect 402102 232938 402186 233174
rect 402422 232938 402454 233174
rect 341794 207218 341826 207454
rect 342062 207218 342146 207454
rect 342382 207218 342414 207454
rect 341794 207134 342414 207218
rect 341794 206898 341826 207134
rect 342062 206898 342146 207134
rect 342382 206898 342414 207134
rect 341794 173454 342414 206898
rect 341794 173218 341826 173454
rect 342062 173218 342146 173454
rect 342382 173218 342414 173454
rect 341794 173134 342414 173218
rect 341794 172898 341826 173134
rect 342062 172898 342146 173134
rect 342382 172898 342414 173134
rect 341794 139454 342414 172898
rect 341794 139218 341826 139454
rect 342062 139218 342146 139454
rect 342382 139218 342414 139454
rect 341794 139134 342414 139218
rect 341794 138898 341826 139134
rect 342062 138898 342146 139134
rect 342382 138898 342414 139134
rect 341794 105454 342414 138898
rect 341794 105218 341826 105454
rect 342062 105218 342146 105454
rect 342382 105218 342414 105454
rect 341794 105134 342414 105218
rect 341794 104898 341826 105134
rect 342062 104898 342146 105134
rect 342382 104898 342414 105134
rect 341794 71454 342414 104898
rect 341794 71218 341826 71454
rect 342062 71218 342146 71454
rect 342382 71218 342414 71454
rect 341794 71134 342414 71218
rect 341794 70898 341826 71134
rect 342062 70898 342146 71134
rect 342382 70898 342414 71134
rect 341794 37454 342414 70898
rect 341794 37218 341826 37454
rect 342062 37218 342146 37454
rect 342382 37218 342414 37454
rect 341794 37134 342414 37218
rect 341794 36898 341826 37134
rect 342062 36898 342146 37134
rect 342382 36898 342414 37134
rect 341794 3454 342414 36898
rect 341794 3218 341826 3454
rect 342062 3218 342146 3454
rect 342382 3218 342414 3454
rect 341794 3134 342414 3218
rect 341794 2898 341826 3134
rect 342062 2898 342146 3134
rect 342382 2898 342414 3134
rect 341794 -346 342414 2898
rect 341794 -582 341826 -346
rect 342062 -582 342146 -346
rect 342382 -582 342414 -346
rect 341794 -666 342414 -582
rect 341794 -902 341826 -666
rect 342062 -902 342146 -666
rect 342382 -902 342414 -666
rect 341794 -7654 342414 -902
rect 345514 211174 346134 214340
rect 345514 210938 345546 211174
rect 345782 210938 345866 211174
rect 346102 210938 346134 211174
rect 345514 210854 346134 210938
rect 345514 210618 345546 210854
rect 345782 210618 345866 210854
rect 346102 210618 346134 210854
rect 345514 177174 346134 210618
rect 345514 176938 345546 177174
rect 345782 176938 345866 177174
rect 346102 176938 346134 177174
rect 345514 176854 346134 176938
rect 345514 176618 345546 176854
rect 345782 176618 345866 176854
rect 346102 176618 346134 176854
rect 345514 143174 346134 176618
rect 345514 142938 345546 143174
rect 345782 142938 345866 143174
rect 346102 142938 346134 143174
rect 345514 142854 346134 142938
rect 345514 142618 345546 142854
rect 345782 142618 345866 142854
rect 346102 142618 346134 142854
rect 345514 109174 346134 142618
rect 345514 108938 345546 109174
rect 345782 108938 345866 109174
rect 346102 108938 346134 109174
rect 345514 108854 346134 108938
rect 345514 108618 345546 108854
rect 345782 108618 345866 108854
rect 346102 108618 346134 108854
rect 345514 75174 346134 108618
rect 345514 74938 345546 75174
rect 345782 74938 345866 75174
rect 346102 74938 346134 75174
rect 345514 74854 346134 74938
rect 345514 74618 345546 74854
rect 345782 74618 345866 74854
rect 346102 74618 346134 74854
rect 345514 41174 346134 74618
rect 345514 40938 345546 41174
rect 345782 40938 345866 41174
rect 346102 40938 346134 41174
rect 345514 40854 346134 40938
rect 345514 40618 345546 40854
rect 345782 40618 345866 40854
rect 346102 40618 346134 40854
rect 345514 7174 346134 40618
rect 345514 6938 345546 7174
rect 345782 6938 345866 7174
rect 346102 6938 346134 7174
rect 345514 6854 346134 6938
rect 345514 6618 345546 6854
rect 345782 6618 345866 6854
rect 346102 6618 346134 6854
rect 345514 -1306 346134 6618
rect 345514 -1542 345546 -1306
rect 345782 -1542 345866 -1306
rect 346102 -1542 346134 -1306
rect 345514 -1626 346134 -1542
rect 345514 -1862 345546 -1626
rect 345782 -1862 345866 -1626
rect 346102 -1862 346134 -1626
rect 345514 -7654 346134 -1862
rect 349234 180894 349854 214340
rect 349234 180658 349266 180894
rect 349502 180658 349586 180894
rect 349822 180658 349854 180894
rect 349234 180574 349854 180658
rect 349234 180338 349266 180574
rect 349502 180338 349586 180574
rect 349822 180338 349854 180574
rect 349234 146894 349854 180338
rect 349234 146658 349266 146894
rect 349502 146658 349586 146894
rect 349822 146658 349854 146894
rect 349234 146574 349854 146658
rect 349234 146338 349266 146574
rect 349502 146338 349586 146574
rect 349822 146338 349854 146574
rect 349234 112894 349854 146338
rect 349234 112658 349266 112894
rect 349502 112658 349586 112894
rect 349822 112658 349854 112894
rect 349234 112574 349854 112658
rect 349234 112338 349266 112574
rect 349502 112338 349586 112574
rect 349822 112338 349854 112574
rect 349234 78894 349854 112338
rect 349234 78658 349266 78894
rect 349502 78658 349586 78894
rect 349822 78658 349854 78894
rect 349234 78574 349854 78658
rect 349234 78338 349266 78574
rect 349502 78338 349586 78574
rect 349822 78338 349854 78574
rect 349234 44894 349854 78338
rect 349234 44658 349266 44894
rect 349502 44658 349586 44894
rect 349822 44658 349854 44894
rect 349234 44574 349854 44658
rect 349234 44338 349266 44574
rect 349502 44338 349586 44574
rect 349822 44338 349854 44574
rect 349234 10894 349854 44338
rect 349234 10658 349266 10894
rect 349502 10658 349586 10894
rect 349822 10658 349854 10894
rect 349234 10574 349854 10658
rect 349234 10338 349266 10574
rect 349502 10338 349586 10574
rect 349822 10338 349854 10574
rect 349234 -2266 349854 10338
rect 349234 -2502 349266 -2266
rect 349502 -2502 349586 -2266
rect 349822 -2502 349854 -2266
rect 349234 -2586 349854 -2502
rect 349234 -2822 349266 -2586
rect 349502 -2822 349586 -2586
rect 349822 -2822 349854 -2586
rect 349234 -7654 349854 -2822
rect 352954 184614 353574 214340
rect 352954 184378 352986 184614
rect 353222 184378 353306 184614
rect 353542 184378 353574 184614
rect 352954 184294 353574 184378
rect 352954 184058 352986 184294
rect 353222 184058 353306 184294
rect 353542 184058 353574 184294
rect 352954 150614 353574 184058
rect 352954 150378 352986 150614
rect 353222 150378 353306 150614
rect 353542 150378 353574 150614
rect 352954 150294 353574 150378
rect 352954 150058 352986 150294
rect 353222 150058 353306 150294
rect 353542 150058 353574 150294
rect 352954 116614 353574 150058
rect 352954 116378 352986 116614
rect 353222 116378 353306 116614
rect 353542 116378 353574 116614
rect 352954 116294 353574 116378
rect 352954 116058 352986 116294
rect 353222 116058 353306 116294
rect 353542 116058 353574 116294
rect 352954 82614 353574 116058
rect 352954 82378 352986 82614
rect 353222 82378 353306 82614
rect 353542 82378 353574 82614
rect 352954 82294 353574 82378
rect 352954 82058 352986 82294
rect 353222 82058 353306 82294
rect 353542 82058 353574 82294
rect 352954 48614 353574 82058
rect 352954 48378 352986 48614
rect 353222 48378 353306 48614
rect 353542 48378 353574 48614
rect 352954 48294 353574 48378
rect 352954 48058 352986 48294
rect 353222 48058 353306 48294
rect 353542 48058 353574 48294
rect 352954 14614 353574 48058
rect 352954 14378 352986 14614
rect 353222 14378 353306 14614
rect 353542 14378 353574 14614
rect 352954 14294 353574 14378
rect 352954 14058 352986 14294
rect 353222 14058 353306 14294
rect 353542 14058 353574 14294
rect 352954 -3226 353574 14058
rect 352954 -3462 352986 -3226
rect 353222 -3462 353306 -3226
rect 353542 -3462 353574 -3226
rect 352954 -3546 353574 -3462
rect 352954 -3782 352986 -3546
rect 353222 -3782 353306 -3546
rect 353542 -3782 353574 -3546
rect 352954 -7654 353574 -3782
rect 356674 188334 357294 214340
rect 356674 188098 356706 188334
rect 356942 188098 357026 188334
rect 357262 188098 357294 188334
rect 356674 188014 357294 188098
rect 356674 187778 356706 188014
rect 356942 187778 357026 188014
rect 357262 187778 357294 188014
rect 356674 154334 357294 187778
rect 356674 154098 356706 154334
rect 356942 154098 357026 154334
rect 357262 154098 357294 154334
rect 356674 154014 357294 154098
rect 356674 153778 356706 154014
rect 356942 153778 357026 154014
rect 357262 153778 357294 154014
rect 356674 120334 357294 153778
rect 356674 120098 356706 120334
rect 356942 120098 357026 120334
rect 357262 120098 357294 120334
rect 356674 120014 357294 120098
rect 356674 119778 356706 120014
rect 356942 119778 357026 120014
rect 357262 119778 357294 120014
rect 356674 86334 357294 119778
rect 356674 86098 356706 86334
rect 356942 86098 357026 86334
rect 357262 86098 357294 86334
rect 356674 86014 357294 86098
rect 356674 85778 356706 86014
rect 356942 85778 357026 86014
rect 357262 85778 357294 86014
rect 356674 52334 357294 85778
rect 356674 52098 356706 52334
rect 356942 52098 357026 52334
rect 357262 52098 357294 52334
rect 356674 52014 357294 52098
rect 356674 51778 356706 52014
rect 356942 51778 357026 52014
rect 357262 51778 357294 52014
rect 356674 18334 357294 51778
rect 356674 18098 356706 18334
rect 356942 18098 357026 18334
rect 357262 18098 357294 18334
rect 356674 18014 357294 18098
rect 356674 17778 356706 18014
rect 356942 17778 357026 18014
rect 357262 17778 357294 18014
rect 356674 -4186 357294 17778
rect 356674 -4422 356706 -4186
rect 356942 -4422 357026 -4186
rect 357262 -4422 357294 -4186
rect 356674 -4506 357294 -4422
rect 356674 -4742 356706 -4506
rect 356942 -4742 357026 -4506
rect 357262 -4742 357294 -4506
rect 356674 -7654 357294 -4742
rect 360394 192054 361014 214340
rect 360394 191818 360426 192054
rect 360662 191818 360746 192054
rect 360982 191818 361014 192054
rect 360394 191734 361014 191818
rect 360394 191498 360426 191734
rect 360662 191498 360746 191734
rect 360982 191498 361014 191734
rect 360394 158054 361014 191498
rect 360394 157818 360426 158054
rect 360662 157818 360746 158054
rect 360982 157818 361014 158054
rect 360394 157734 361014 157818
rect 360394 157498 360426 157734
rect 360662 157498 360746 157734
rect 360982 157498 361014 157734
rect 360394 124054 361014 157498
rect 360394 123818 360426 124054
rect 360662 123818 360746 124054
rect 360982 123818 361014 124054
rect 360394 123734 361014 123818
rect 360394 123498 360426 123734
rect 360662 123498 360746 123734
rect 360982 123498 361014 123734
rect 360394 90054 361014 123498
rect 360394 89818 360426 90054
rect 360662 89818 360746 90054
rect 360982 89818 361014 90054
rect 360394 89734 361014 89818
rect 360394 89498 360426 89734
rect 360662 89498 360746 89734
rect 360982 89498 361014 89734
rect 360394 56054 361014 89498
rect 360394 55818 360426 56054
rect 360662 55818 360746 56054
rect 360982 55818 361014 56054
rect 360394 55734 361014 55818
rect 360394 55498 360426 55734
rect 360662 55498 360746 55734
rect 360982 55498 361014 55734
rect 360394 22054 361014 55498
rect 360394 21818 360426 22054
rect 360662 21818 360746 22054
rect 360982 21818 361014 22054
rect 360394 21734 361014 21818
rect 360394 21498 360426 21734
rect 360662 21498 360746 21734
rect 360982 21498 361014 21734
rect 360394 -5146 361014 21498
rect 360394 -5382 360426 -5146
rect 360662 -5382 360746 -5146
rect 360982 -5382 361014 -5146
rect 360394 -5466 361014 -5382
rect 360394 -5702 360426 -5466
rect 360662 -5702 360746 -5466
rect 360982 -5702 361014 -5466
rect 360394 -7654 361014 -5702
rect 364114 195774 364734 214340
rect 364114 195538 364146 195774
rect 364382 195538 364466 195774
rect 364702 195538 364734 195774
rect 364114 195454 364734 195538
rect 364114 195218 364146 195454
rect 364382 195218 364466 195454
rect 364702 195218 364734 195454
rect 364114 161774 364734 195218
rect 364114 161538 364146 161774
rect 364382 161538 364466 161774
rect 364702 161538 364734 161774
rect 364114 161454 364734 161538
rect 364114 161218 364146 161454
rect 364382 161218 364466 161454
rect 364702 161218 364734 161454
rect 364114 127774 364734 161218
rect 364114 127538 364146 127774
rect 364382 127538 364466 127774
rect 364702 127538 364734 127774
rect 364114 127454 364734 127538
rect 364114 127218 364146 127454
rect 364382 127218 364466 127454
rect 364702 127218 364734 127454
rect 364114 93774 364734 127218
rect 364114 93538 364146 93774
rect 364382 93538 364466 93774
rect 364702 93538 364734 93774
rect 364114 93454 364734 93538
rect 364114 93218 364146 93454
rect 364382 93218 364466 93454
rect 364702 93218 364734 93454
rect 364114 59774 364734 93218
rect 364114 59538 364146 59774
rect 364382 59538 364466 59774
rect 364702 59538 364734 59774
rect 364114 59454 364734 59538
rect 364114 59218 364146 59454
rect 364382 59218 364466 59454
rect 364702 59218 364734 59454
rect 364114 25774 364734 59218
rect 364114 25538 364146 25774
rect 364382 25538 364466 25774
rect 364702 25538 364734 25774
rect 364114 25454 364734 25538
rect 364114 25218 364146 25454
rect 364382 25218 364466 25454
rect 364702 25218 364734 25454
rect 364114 -6106 364734 25218
rect 364114 -6342 364146 -6106
rect 364382 -6342 364466 -6106
rect 364702 -6342 364734 -6106
rect 364114 -6426 364734 -6342
rect 364114 -6662 364146 -6426
rect 364382 -6662 364466 -6426
rect 364702 -6662 364734 -6426
rect 364114 -7654 364734 -6662
rect 367834 199494 368454 214340
rect 367834 199258 367866 199494
rect 368102 199258 368186 199494
rect 368422 199258 368454 199494
rect 367834 199174 368454 199258
rect 367834 198938 367866 199174
rect 368102 198938 368186 199174
rect 368422 198938 368454 199174
rect 367834 165494 368454 198938
rect 367834 165258 367866 165494
rect 368102 165258 368186 165494
rect 368422 165258 368454 165494
rect 367834 165174 368454 165258
rect 367834 164938 367866 165174
rect 368102 164938 368186 165174
rect 368422 164938 368454 165174
rect 367834 131494 368454 164938
rect 367834 131258 367866 131494
rect 368102 131258 368186 131494
rect 368422 131258 368454 131494
rect 367834 131174 368454 131258
rect 367834 130938 367866 131174
rect 368102 130938 368186 131174
rect 368422 130938 368454 131174
rect 367834 97494 368454 130938
rect 367834 97258 367866 97494
rect 368102 97258 368186 97494
rect 368422 97258 368454 97494
rect 367834 97174 368454 97258
rect 367834 96938 367866 97174
rect 368102 96938 368186 97174
rect 368422 96938 368454 97174
rect 367834 63494 368454 96938
rect 367834 63258 367866 63494
rect 368102 63258 368186 63494
rect 368422 63258 368454 63494
rect 367834 63174 368454 63258
rect 367834 62938 367866 63174
rect 368102 62938 368186 63174
rect 368422 62938 368454 63174
rect 367834 29494 368454 62938
rect 367834 29258 367866 29494
rect 368102 29258 368186 29494
rect 368422 29258 368454 29494
rect 367834 29174 368454 29258
rect 367834 28938 367866 29174
rect 368102 28938 368186 29174
rect 368422 28938 368454 29174
rect 367834 -7066 368454 28938
rect 367834 -7302 367866 -7066
rect 368102 -7302 368186 -7066
rect 368422 -7302 368454 -7066
rect 367834 -7386 368454 -7302
rect 367834 -7622 367866 -7386
rect 368102 -7622 368186 -7386
rect 368422 -7622 368454 -7386
rect 367834 -7654 368454 -7622
rect 375794 207454 376414 214340
rect 375794 207218 375826 207454
rect 376062 207218 376146 207454
rect 376382 207218 376414 207454
rect 375794 207134 376414 207218
rect 375794 206898 375826 207134
rect 376062 206898 376146 207134
rect 376382 206898 376414 207134
rect 375794 173454 376414 206898
rect 375794 173218 375826 173454
rect 376062 173218 376146 173454
rect 376382 173218 376414 173454
rect 375794 173134 376414 173218
rect 375794 172898 375826 173134
rect 376062 172898 376146 173134
rect 376382 172898 376414 173134
rect 375794 139454 376414 172898
rect 375794 139218 375826 139454
rect 376062 139218 376146 139454
rect 376382 139218 376414 139454
rect 375794 139134 376414 139218
rect 375794 138898 375826 139134
rect 376062 138898 376146 139134
rect 376382 138898 376414 139134
rect 375794 105454 376414 138898
rect 375794 105218 375826 105454
rect 376062 105218 376146 105454
rect 376382 105218 376414 105454
rect 375794 105134 376414 105218
rect 375794 104898 375826 105134
rect 376062 104898 376146 105134
rect 376382 104898 376414 105134
rect 375794 71454 376414 104898
rect 375794 71218 375826 71454
rect 376062 71218 376146 71454
rect 376382 71218 376414 71454
rect 375794 71134 376414 71218
rect 375794 70898 375826 71134
rect 376062 70898 376146 71134
rect 376382 70898 376414 71134
rect 375794 37454 376414 70898
rect 375794 37218 375826 37454
rect 376062 37218 376146 37454
rect 376382 37218 376414 37454
rect 375794 37134 376414 37218
rect 375794 36898 375826 37134
rect 376062 36898 376146 37134
rect 376382 36898 376414 37134
rect 375794 3454 376414 36898
rect 375794 3218 375826 3454
rect 376062 3218 376146 3454
rect 376382 3218 376414 3454
rect 375794 3134 376414 3218
rect 375794 2898 375826 3134
rect 376062 2898 376146 3134
rect 376382 2898 376414 3134
rect 375794 -346 376414 2898
rect 375794 -582 375826 -346
rect 376062 -582 376146 -346
rect 376382 -582 376414 -346
rect 375794 -666 376414 -582
rect 375794 -902 375826 -666
rect 376062 -902 376146 -666
rect 376382 -902 376414 -666
rect 375794 -7654 376414 -902
rect 379514 211174 380134 214340
rect 379514 210938 379546 211174
rect 379782 210938 379866 211174
rect 380102 210938 380134 211174
rect 379514 210854 380134 210938
rect 379514 210618 379546 210854
rect 379782 210618 379866 210854
rect 380102 210618 380134 210854
rect 379514 177174 380134 210618
rect 379514 176938 379546 177174
rect 379782 176938 379866 177174
rect 380102 176938 380134 177174
rect 379514 176854 380134 176938
rect 379514 176618 379546 176854
rect 379782 176618 379866 176854
rect 380102 176618 380134 176854
rect 379514 143174 380134 176618
rect 379514 142938 379546 143174
rect 379782 142938 379866 143174
rect 380102 142938 380134 143174
rect 379514 142854 380134 142938
rect 379514 142618 379546 142854
rect 379782 142618 379866 142854
rect 380102 142618 380134 142854
rect 379514 109174 380134 142618
rect 379514 108938 379546 109174
rect 379782 108938 379866 109174
rect 380102 108938 380134 109174
rect 379514 108854 380134 108938
rect 379514 108618 379546 108854
rect 379782 108618 379866 108854
rect 380102 108618 380134 108854
rect 379514 75174 380134 108618
rect 379514 74938 379546 75174
rect 379782 74938 379866 75174
rect 380102 74938 380134 75174
rect 379514 74854 380134 74938
rect 379514 74618 379546 74854
rect 379782 74618 379866 74854
rect 380102 74618 380134 74854
rect 379514 41174 380134 74618
rect 379514 40938 379546 41174
rect 379782 40938 379866 41174
rect 380102 40938 380134 41174
rect 379514 40854 380134 40938
rect 379514 40618 379546 40854
rect 379782 40618 379866 40854
rect 380102 40618 380134 40854
rect 379514 7174 380134 40618
rect 379514 6938 379546 7174
rect 379782 6938 379866 7174
rect 380102 6938 380134 7174
rect 379514 6854 380134 6938
rect 379514 6618 379546 6854
rect 379782 6618 379866 6854
rect 380102 6618 380134 6854
rect 379514 -1306 380134 6618
rect 379514 -1542 379546 -1306
rect 379782 -1542 379866 -1306
rect 380102 -1542 380134 -1306
rect 379514 -1626 380134 -1542
rect 379514 -1862 379546 -1626
rect 379782 -1862 379866 -1626
rect 380102 -1862 380134 -1626
rect 379514 -7654 380134 -1862
rect 383234 180894 383854 214340
rect 383234 180658 383266 180894
rect 383502 180658 383586 180894
rect 383822 180658 383854 180894
rect 383234 180574 383854 180658
rect 383234 180338 383266 180574
rect 383502 180338 383586 180574
rect 383822 180338 383854 180574
rect 383234 146894 383854 180338
rect 383234 146658 383266 146894
rect 383502 146658 383586 146894
rect 383822 146658 383854 146894
rect 383234 146574 383854 146658
rect 383234 146338 383266 146574
rect 383502 146338 383586 146574
rect 383822 146338 383854 146574
rect 383234 112894 383854 146338
rect 383234 112658 383266 112894
rect 383502 112658 383586 112894
rect 383822 112658 383854 112894
rect 383234 112574 383854 112658
rect 383234 112338 383266 112574
rect 383502 112338 383586 112574
rect 383822 112338 383854 112574
rect 383234 78894 383854 112338
rect 383234 78658 383266 78894
rect 383502 78658 383586 78894
rect 383822 78658 383854 78894
rect 383234 78574 383854 78658
rect 383234 78338 383266 78574
rect 383502 78338 383586 78574
rect 383822 78338 383854 78574
rect 383234 44894 383854 78338
rect 383234 44658 383266 44894
rect 383502 44658 383586 44894
rect 383822 44658 383854 44894
rect 383234 44574 383854 44658
rect 383234 44338 383266 44574
rect 383502 44338 383586 44574
rect 383822 44338 383854 44574
rect 383234 10894 383854 44338
rect 383234 10658 383266 10894
rect 383502 10658 383586 10894
rect 383822 10658 383854 10894
rect 383234 10574 383854 10658
rect 383234 10338 383266 10574
rect 383502 10338 383586 10574
rect 383822 10338 383854 10574
rect 383234 -2266 383854 10338
rect 383234 -2502 383266 -2266
rect 383502 -2502 383586 -2266
rect 383822 -2502 383854 -2266
rect 383234 -2586 383854 -2502
rect 383234 -2822 383266 -2586
rect 383502 -2822 383586 -2586
rect 383822 -2822 383854 -2586
rect 383234 -7654 383854 -2822
rect 386954 184614 387574 214340
rect 386954 184378 386986 184614
rect 387222 184378 387306 184614
rect 387542 184378 387574 184614
rect 386954 184294 387574 184378
rect 386954 184058 386986 184294
rect 387222 184058 387306 184294
rect 387542 184058 387574 184294
rect 386954 150614 387574 184058
rect 386954 150378 386986 150614
rect 387222 150378 387306 150614
rect 387542 150378 387574 150614
rect 386954 150294 387574 150378
rect 386954 150058 386986 150294
rect 387222 150058 387306 150294
rect 387542 150058 387574 150294
rect 386954 116614 387574 150058
rect 386954 116378 386986 116614
rect 387222 116378 387306 116614
rect 387542 116378 387574 116614
rect 386954 116294 387574 116378
rect 386954 116058 386986 116294
rect 387222 116058 387306 116294
rect 387542 116058 387574 116294
rect 386954 82614 387574 116058
rect 386954 82378 386986 82614
rect 387222 82378 387306 82614
rect 387542 82378 387574 82614
rect 386954 82294 387574 82378
rect 386954 82058 386986 82294
rect 387222 82058 387306 82294
rect 387542 82058 387574 82294
rect 386954 48614 387574 82058
rect 386954 48378 386986 48614
rect 387222 48378 387306 48614
rect 387542 48378 387574 48614
rect 386954 48294 387574 48378
rect 386954 48058 386986 48294
rect 387222 48058 387306 48294
rect 387542 48058 387574 48294
rect 386954 14614 387574 48058
rect 386954 14378 386986 14614
rect 387222 14378 387306 14614
rect 387542 14378 387574 14614
rect 386954 14294 387574 14378
rect 386954 14058 386986 14294
rect 387222 14058 387306 14294
rect 387542 14058 387574 14294
rect 386954 -3226 387574 14058
rect 386954 -3462 386986 -3226
rect 387222 -3462 387306 -3226
rect 387542 -3462 387574 -3226
rect 386954 -3546 387574 -3462
rect 386954 -3782 386986 -3546
rect 387222 -3782 387306 -3546
rect 387542 -3782 387574 -3546
rect 386954 -7654 387574 -3782
rect 390674 188334 391294 214340
rect 390674 188098 390706 188334
rect 390942 188098 391026 188334
rect 391262 188098 391294 188334
rect 390674 188014 391294 188098
rect 390674 187778 390706 188014
rect 390942 187778 391026 188014
rect 391262 187778 391294 188014
rect 390674 154334 391294 187778
rect 390674 154098 390706 154334
rect 390942 154098 391026 154334
rect 391262 154098 391294 154334
rect 390674 154014 391294 154098
rect 390674 153778 390706 154014
rect 390942 153778 391026 154014
rect 391262 153778 391294 154014
rect 390674 120334 391294 153778
rect 390674 120098 390706 120334
rect 390942 120098 391026 120334
rect 391262 120098 391294 120334
rect 390674 120014 391294 120098
rect 390674 119778 390706 120014
rect 390942 119778 391026 120014
rect 391262 119778 391294 120014
rect 390674 86334 391294 119778
rect 390674 86098 390706 86334
rect 390942 86098 391026 86334
rect 391262 86098 391294 86334
rect 390674 86014 391294 86098
rect 390674 85778 390706 86014
rect 390942 85778 391026 86014
rect 391262 85778 391294 86014
rect 390674 52334 391294 85778
rect 390674 52098 390706 52334
rect 390942 52098 391026 52334
rect 391262 52098 391294 52334
rect 390674 52014 391294 52098
rect 390674 51778 390706 52014
rect 390942 51778 391026 52014
rect 391262 51778 391294 52014
rect 390674 18334 391294 51778
rect 390674 18098 390706 18334
rect 390942 18098 391026 18334
rect 391262 18098 391294 18334
rect 390674 18014 391294 18098
rect 390674 17778 390706 18014
rect 390942 17778 391026 18014
rect 391262 17778 391294 18014
rect 390674 -4186 391294 17778
rect 390674 -4422 390706 -4186
rect 390942 -4422 391026 -4186
rect 391262 -4422 391294 -4186
rect 390674 -4506 391294 -4422
rect 390674 -4742 390706 -4506
rect 390942 -4742 391026 -4506
rect 391262 -4742 391294 -4506
rect 390674 -7654 391294 -4742
rect 394394 192054 395014 214340
rect 394394 191818 394426 192054
rect 394662 191818 394746 192054
rect 394982 191818 395014 192054
rect 394394 191734 395014 191818
rect 394394 191498 394426 191734
rect 394662 191498 394746 191734
rect 394982 191498 395014 191734
rect 394394 158054 395014 191498
rect 394394 157818 394426 158054
rect 394662 157818 394746 158054
rect 394982 157818 395014 158054
rect 394394 157734 395014 157818
rect 394394 157498 394426 157734
rect 394662 157498 394746 157734
rect 394982 157498 395014 157734
rect 394394 124054 395014 157498
rect 394394 123818 394426 124054
rect 394662 123818 394746 124054
rect 394982 123818 395014 124054
rect 394394 123734 395014 123818
rect 394394 123498 394426 123734
rect 394662 123498 394746 123734
rect 394982 123498 395014 123734
rect 394394 90054 395014 123498
rect 394394 89818 394426 90054
rect 394662 89818 394746 90054
rect 394982 89818 395014 90054
rect 394394 89734 395014 89818
rect 394394 89498 394426 89734
rect 394662 89498 394746 89734
rect 394982 89498 395014 89734
rect 394394 56054 395014 89498
rect 394394 55818 394426 56054
rect 394662 55818 394746 56054
rect 394982 55818 395014 56054
rect 394394 55734 395014 55818
rect 394394 55498 394426 55734
rect 394662 55498 394746 55734
rect 394982 55498 395014 55734
rect 394394 22054 395014 55498
rect 394394 21818 394426 22054
rect 394662 21818 394746 22054
rect 394982 21818 395014 22054
rect 394394 21734 395014 21818
rect 394394 21498 394426 21734
rect 394662 21498 394746 21734
rect 394982 21498 395014 21734
rect 394394 -5146 395014 21498
rect 394394 -5382 394426 -5146
rect 394662 -5382 394746 -5146
rect 394982 -5382 395014 -5146
rect 394394 -5466 395014 -5382
rect 394394 -5702 394426 -5466
rect 394662 -5702 394746 -5466
rect 394982 -5702 395014 -5466
rect 394394 -7654 395014 -5702
rect 398114 195774 398734 214340
rect 398114 195538 398146 195774
rect 398382 195538 398466 195774
rect 398702 195538 398734 195774
rect 398114 195454 398734 195538
rect 398114 195218 398146 195454
rect 398382 195218 398466 195454
rect 398702 195218 398734 195454
rect 398114 161774 398734 195218
rect 398114 161538 398146 161774
rect 398382 161538 398466 161774
rect 398702 161538 398734 161774
rect 398114 161454 398734 161538
rect 398114 161218 398146 161454
rect 398382 161218 398466 161454
rect 398702 161218 398734 161454
rect 398114 127774 398734 161218
rect 398114 127538 398146 127774
rect 398382 127538 398466 127774
rect 398702 127538 398734 127774
rect 398114 127454 398734 127538
rect 398114 127218 398146 127454
rect 398382 127218 398466 127454
rect 398702 127218 398734 127454
rect 398114 93774 398734 127218
rect 398114 93538 398146 93774
rect 398382 93538 398466 93774
rect 398702 93538 398734 93774
rect 398114 93454 398734 93538
rect 398114 93218 398146 93454
rect 398382 93218 398466 93454
rect 398702 93218 398734 93454
rect 398114 59774 398734 93218
rect 398114 59538 398146 59774
rect 398382 59538 398466 59774
rect 398702 59538 398734 59774
rect 398114 59454 398734 59538
rect 398114 59218 398146 59454
rect 398382 59218 398466 59454
rect 398702 59218 398734 59454
rect 398114 25774 398734 59218
rect 398114 25538 398146 25774
rect 398382 25538 398466 25774
rect 398702 25538 398734 25774
rect 398114 25454 398734 25538
rect 398114 25218 398146 25454
rect 398382 25218 398466 25454
rect 398702 25218 398734 25454
rect 398114 -6106 398734 25218
rect 398114 -6342 398146 -6106
rect 398382 -6342 398466 -6106
rect 398702 -6342 398734 -6106
rect 398114 -6426 398734 -6342
rect 398114 -6662 398146 -6426
rect 398382 -6662 398466 -6426
rect 398702 -6662 398734 -6426
rect 398114 -7654 398734 -6662
rect 401834 199494 402454 232938
rect 401834 199258 401866 199494
rect 402102 199258 402186 199494
rect 402422 199258 402454 199494
rect 401834 199174 402454 199258
rect 401834 198938 401866 199174
rect 402102 198938 402186 199174
rect 402422 198938 402454 199174
rect 401834 165494 402454 198938
rect 401834 165258 401866 165494
rect 402102 165258 402186 165494
rect 402422 165258 402454 165494
rect 401834 165174 402454 165258
rect 401834 164938 401866 165174
rect 402102 164938 402186 165174
rect 402422 164938 402454 165174
rect 401834 131494 402454 164938
rect 401834 131258 401866 131494
rect 402102 131258 402186 131494
rect 402422 131258 402454 131494
rect 401834 131174 402454 131258
rect 401834 130938 401866 131174
rect 402102 130938 402186 131174
rect 402422 130938 402454 131174
rect 401834 97494 402454 130938
rect 401834 97258 401866 97494
rect 402102 97258 402186 97494
rect 402422 97258 402454 97494
rect 401834 97174 402454 97258
rect 401834 96938 401866 97174
rect 402102 96938 402186 97174
rect 402422 96938 402454 97174
rect 401834 63494 402454 96938
rect 401834 63258 401866 63494
rect 402102 63258 402186 63494
rect 402422 63258 402454 63494
rect 401834 63174 402454 63258
rect 401834 62938 401866 63174
rect 402102 62938 402186 63174
rect 402422 62938 402454 63174
rect 401834 29494 402454 62938
rect 401834 29258 401866 29494
rect 402102 29258 402186 29494
rect 402422 29258 402454 29494
rect 401834 29174 402454 29258
rect 401834 28938 401866 29174
rect 402102 28938 402186 29174
rect 402422 28938 402454 29174
rect 401834 -7066 402454 28938
rect 401834 -7302 401866 -7066
rect 402102 -7302 402186 -7066
rect 402422 -7302 402454 -7066
rect 401834 -7386 402454 -7302
rect 401834 -7622 401866 -7386
rect 402102 -7622 402186 -7386
rect 402422 -7622 402454 -7386
rect 401834 -7654 402454 -7622
rect 409794 704838 410414 711590
rect 409794 704602 409826 704838
rect 410062 704602 410146 704838
rect 410382 704602 410414 704838
rect 409794 704518 410414 704602
rect 409794 704282 409826 704518
rect 410062 704282 410146 704518
rect 410382 704282 410414 704518
rect 409794 683454 410414 704282
rect 409794 683218 409826 683454
rect 410062 683218 410146 683454
rect 410382 683218 410414 683454
rect 409794 683134 410414 683218
rect 409794 682898 409826 683134
rect 410062 682898 410146 683134
rect 410382 682898 410414 683134
rect 409794 649454 410414 682898
rect 409794 649218 409826 649454
rect 410062 649218 410146 649454
rect 410382 649218 410414 649454
rect 409794 649134 410414 649218
rect 409794 648898 409826 649134
rect 410062 648898 410146 649134
rect 410382 648898 410414 649134
rect 409794 615454 410414 648898
rect 409794 615218 409826 615454
rect 410062 615218 410146 615454
rect 410382 615218 410414 615454
rect 409794 615134 410414 615218
rect 409794 614898 409826 615134
rect 410062 614898 410146 615134
rect 410382 614898 410414 615134
rect 409794 581454 410414 614898
rect 409794 581218 409826 581454
rect 410062 581218 410146 581454
rect 410382 581218 410414 581454
rect 409794 581134 410414 581218
rect 409794 580898 409826 581134
rect 410062 580898 410146 581134
rect 410382 580898 410414 581134
rect 409794 547454 410414 580898
rect 409794 547218 409826 547454
rect 410062 547218 410146 547454
rect 410382 547218 410414 547454
rect 409794 547134 410414 547218
rect 409794 546898 409826 547134
rect 410062 546898 410146 547134
rect 410382 546898 410414 547134
rect 409794 513454 410414 546898
rect 409794 513218 409826 513454
rect 410062 513218 410146 513454
rect 410382 513218 410414 513454
rect 409794 513134 410414 513218
rect 409794 512898 409826 513134
rect 410062 512898 410146 513134
rect 410382 512898 410414 513134
rect 409794 479454 410414 512898
rect 409794 479218 409826 479454
rect 410062 479218 410146 479454
rect 410382 479218 410414 479454
rect 409794 479134 410414 479218
rect 409794 478898 409826 479134
rect 410062 478898 410146 479134
rect 410382 478898 410414 479134
rect 409794 445454 410414 478898
rect 409794 445218 409826 445454
rect 410062 445218 410146 445454
rect 410382 445218 410414 445454
rect 409794 445134 410414 445218
rect 409794 444898 409826 445134
rect 410062 444898 410146 445134
rect 410382 444898 410414 445134
rect 409794 411454 410414 444898
rect 409794 411218 409826 411454
rect 410062 411218 410146 411454
rect 410382 411218 410414 411454
rect 409794 411134 410414 411218
rect 409794 410898 409826 411134
rect 410062 410898 410146 411134
rect 410382 410898 410414 411134
rect 409794 377454 410414 410898
rect 409794 377218 409826 377454
rect 410062 377218 410146 377454
rect 410382 377218 410414 377454
rect 409794 377134 410414 377218
rect 409794 376898 409826 377134
rect 410062 376898 410146 377134
rect 410382 376898 410414 377134
rect 409794 343454 410414 376898
rect 409794 343218 409826 343454
rect 410062 343218 410146 343454
rect 410382 343218 410414 343454
rect 409794 343134 410414 343218
rect 409794 342898 409826 343134
rect 410062 342898 410146 343134
rect 410382 342898 410414 343134
rect 409794 309454 410414 342898
rect 409794 309218 409826 309454
rect 410062 309218 410146 309454
rect 410382 309218 410414 309454
rect 409794 309134 410414 309218
rect 409794 308898 409826 309134
rect 410062 308898 410146 309134
rect 410382 308898 410414 309134
rect 409794 275454 410414 308898
rect 409794 275218 409826 275454
rect 410062 275218 410146 275454
rect 410382 275218 410414 275454
rect 409794 275134 410414 275218
rect 409794 274898 409826 275134
rect 410062 274898 410146 275134
rect 410382 274898 410414 275134
rect 409794 241454 410414 274898
rect 409794 241218 409826 241454
rect 410062 241218 410146 241454
rect 410382 241218 410414 241454
rect 409794 241134 410414 241218
rect 409794 240898 409826 241134
rect 410062 240898 410146 241134
rect 410382 240898 410414 241134
rect 409794 207454 410414 240898
rect 409794 207218 409826 207454
rect 410062 207218 410146 207454
rect 410382 207218 410414 207454
rect 409794 207134 410414 207218
rect 409794 206898 409826 207134
rect 410062 206898 410146 207134
rect 410382 206898 410414 207134
rect 409794 173454 410414 206898
rect 409794 173218 409826 173454
rect 410062 173218 410146 173454
rect 410382 173218 410414 173454
rect 409794 173134 410414 173218
rect 409794 172898 409826 173134
rect 410062 172898 410146 173134
rect 410382 172898 410414 173134
rect 409794 139454 410414 172898
rect 409794 139218 409826 139454
rect 410062 139218 410146 139454
rect 410382 139218 410414 139454
rect 409794 139134 410414 139218
rect 409794 138898 409826 139134
rect 410062 138898 410146 139134
rect 410382 138898 410414 139134
rect 409794 105454 410414 138898
rect 409794 105218 409826 105454
rect 410062 105218 410146 105454
rect 410382 105218 410414 105454
rect 409794 105134 410414 105218
rect 409794 104898 409826 105134
rect 410062 104898 410146 105134
rect 410382 104898 410414 105134
rect 409794 71454 410414 104898
rect 409794 71218 409826 71454
rect 410062 71218 410146 71454
rect 410382 71218 410414 71454
rect 409794 71134 410414 71218
rect 409794 70898 409826 71134
rect 410062 70898 410146 71134
rect 410382 70898 410414 71134
rect 409794 37454 410414 70898
rect 409794 37218 409826 37454
rect 410062 37218 410146 37454
rect 410382 37218 410414 37454
rect 409794 37134 410414 37218
rect 409794 36898 409826 37134
rect 410062 36898 410146 37134
rect 410382 36898 410414 37134
rect 409794 3454 410414 36898
rect 409794 3218 409826 3454
rect 410062 3218 410146 3454
rect 410382 3218 410414 3454
rect 409794 3134 410414 3218
rect 409794 2898 409826 3134
rect 410062 2898 410146 3134
rect 410382 2898 410414 3134
rect 409794 -346 410414 2898
rect 409794 -582 409826 -346
rect 410062 -582 410146 -346
rect 410382 -582 410414 -346
rect 409794 -666 410414 -582
rect 409794 -902 409826 -666
rect 410062 -902 410146 -666
rect 410382 -902 410414 -666
rect 409794 -7654 410414 -902
rect 413514 705798 414134 711590
rect 413514 705562 413546 705798
rect 413782 705562 413866 705798
rect 414102 705562 414134 705798
rect 413514 705478 414134 705562
rect 413514 705242 413546 705478
rect 413782 705242 413866 705478
rect 414102 705242 414134 705478
rect 413514 687174 414134 705242
rect 413514 686938 413546 687174
rect 413782 686938 413866 687174
rect 414102 686938 414134 687174
rect 413514 686854 414134 686938
rect 413514 686618 413546 686854
rect 413782 686618 413866 686854
rect 414102 686618 414134 686854
rect 413514 653174 414134 686618
rect 413514 652938 413546 653174
rect 413782 652938 413866 653174
rect 414102 652938 414134 653174
rect 413514 652854 414134 652938
rect 413514 652618 413546 652854
rect 413782 652618 413866 652854
rect 414102 652618 414134 652854
rect 413514 619174 414134 652618
rect 413514 618938 413546 619174
rect 413782 618938 413866 619174
rect 414102 618938 414134 619174
rect 413514 618854 414134 618938
rect 413514 618618 413546 618854
rect 413782 618618 413866 618854
rect 414102 618618 414134 618854
rect 413514 585174 414134 618618
rect 413514 584938 413546 585174
rect 413782 584938 413866 585174
rect 414102 584938 414134 585174
rect 413514 584854 414134 584938
rect 413514 584618 413546 584854
rect 413782 584618 413866 584854
rect 414102 584618 414134 584854
rect 413514 551174 414134 584618
rect 413514 550938 413546 551174
rect 413782 550938 413866 551174
rect 414102 550938 414134 551174
rect 413514 550854 414134 550938
rect 413514 550618 413546 550854
rect 413782 550618 413866 550854
rect 414102 550618 414134 550854
rect 413514 517174 414134 550618
rect 413514 516938 413546 517174
rect 413782 516938 413866 517174
rect 414102 516938 414134 517174
rect 413514 516854 414134 516938
rect 413514 516618 413546 516854
rect 413782 516618 413866 516854
rect 414102 516618 414134 516854
rect 413514 483174 414134 516618
rect 413514 482938 413546 483174
rect 413782 482938 413866 483174
rect 414102 482938 414134 483174
rect 413514 482854 414134 482938
rect 413514 482618 413546 482854
rect 413782 482618 413866 482854
rect 414102 482618 414134 482854
rect 413514 449174 414134 482618
rect 413514 448938 413546 449174
rect 413782 448938 413866 449174
rect 414102 448938 414134 449174
rect 413514 448854 414134 448938
rect 413514 448618 413546 448854
rect 413782 448618 413866 448854
rect 414102 448618 414134 448854
rect 413514 415174 414134 448618
rect 413514 414938 413546 415174
rect 413782 414938 413866 415174
rect 414102 414938 414134 415174
rect 413514 414854 414134 414938
rect 413514 414618 413546 414854
rect 413782 414618 413866 414854
rect 414102 414618 414134 414854
rect 413514 381174 414134 414618
rect 413514 380938 413546 381174
rect 413782 380938 413866 381174
rect 414102 380938 414134 381174
rect 413514 380854 414134 380938
rect 413514 380618 413546 380854
rect 413782 380618 413866 380854
rect 414102 380618 414134 380854
rect 413514 347174 414134 380618
rect 413514 346938 413546 347174
rect 413782 346938 413866 347174
rect 414102 346938 414134 347174
rect 413514 346854 414134 346938
rect 413514 346618 413546 346854
rect 413782 346618 413866 346854
rect 414102 346618 414134 346854
rect 413514 313174 414134 346618
rect 413514 312938 413546 313174
rect 413782 312938 413866 313174
rect 414102 312938 414134 313174
rect 413514 312854 414134 312938
rect 413514 312618 413546 312854
rect 413782 312618 413866 312854
rect 414102 312618 414134 312854
rect 413514 279174 414134 312618
rect 413514 278938 413546 279174
rect 413782 278938 413866 279174
rect 414102 278938 414134 279174
rect 413514 278854 414134 278938
rect 413514 278618 413546 278854
rect 413782 278618 413866 278854
rect 414102 278618 414134 278854
rect 413514 245174 414134 278618
rect 413514 244938 413546 245174
rect 413782 244938 413866 245174
rect 414102 244938 414134 245174
rect 413514 244854 414134 244938
rect 413514 244618 413546 244854
rect 413782 244618 413866 244854
rect 414102 244618 414134 244854
rect 413514 211174 414134 244618
rect 413514 210938 413546 211174
rect 413782 210938 413866 211174
rect 414102 210938 414134 211174
rect 413514 210854 414134 210938
rect 413514 210618 413546 210854
rect 413782 210618 413866 210854
rect 414102 210618 414134 210854
rect 413514 177174 414134 210618
rect 413514 176938 413546 177174
rect 413782 176938 413866 177174
rect 414102 176938 414134 177174
rect 413514 176854 414134 176938
rect 413514 176618 413546 176854
rect 413782 176618 413866 176854
rect 414102 176618 414134 176854
rect 413514 143174 414134 176618
rect 413514 142938 413546 143174
rect 413782 142938 413866 143174
rect 414102 142938 414134 143174
rect 413514 142854 414134 142938
rect 413514 142618 413546 142854
rect 413782 142618 413866 142854
rect 414102 142618 414134 142854
rect 413514 109174 414134 142618
rect 413514 108938 413546 109174
rect 413782 108938 413866 109174
rect 414102 108938 414134 109174
rect 413514 108854 414134 108938
rect 413514 108618 413546 108854
rect 413782 108618 413866 108854
rect 414102 108618 414134 108854
rect 413514 75174 414134 108618
rect 413514 74938 413546 75174
rect 413782 74938 413866 75174
rect 414102 74938 414134 75174
rect 413514 74854 414134 74938
rect 413514 74618 413546 74854
rect 413782 74618 413866 74854
rect 414102 74618 414134 74854
rect 413514 41174 414134 74618
rect 413514 40938 413546 41174
rect 413782 40938 413866 41174
rect 414102 40938 414134 41174
rect 413514 40854 414134 40938
rect 413514 40618 413546 40854
rect 413782 40618 413866 40854
rect 414102 40618 414134 40854
rect 413514 7174 414134 40618
rect 413514 6938 413546 7174
rect 413782 6938 413866 7174
rect 414102 6938 414134 7174
rect 413514 6854 414134 6938
rect 413514 6618 413546 6854
rect 413782 6618 413866 6854
rect 414102 6618 414134 6854
rect 413514 -1306 414134 6618
rect 413514 -1542 413546 -1306
rect 413782 -1542 413866 -1306
rect 414102 -1542 414134 -1306
rect 413514 -1626 414134 -1542
rect 413514 -1862 413546 -1626
rect 413782 -1862 413866 -1626
rect 414102 -1862 414134 -1626
rect 413514 -7654 414134 -1862
rect 417234 706758 417854 711590
rect 417234 706522 417266 706758
rect 417502 706522 417586 706758
rect 417822 706522 417854 706758
rect 417234 706438 417854 706522
rect 417234 706202 417266 706438
rect 417502 706202 417586 706438
rect 417822 706202 417854 706438
rect 417234 690894 417854 706202
rect 417234 690658 417266 690894
rect 417502 690658 417586 690894
rect 417822 690658 417854 690894
rect 417234 690574 417854 690658
rect 417234 690338 417266 690574
rect 417502 690338 417586 690574
rect 417822 690338 417854 690574
rect 417234 656894 417854 690338
rect 417234 656658 417266 656894
rect 417502 656658 417586 656894
rect 417822 656658 417854 656894
rect 417234 656574 417854 656658
rect 417234 656338 417266 656574
rect 417502 656338 417586 656574
rect 417822 656338 417854 656574
rect 417234 622894 417854 656338
rect 417234 622658 417266 622894
rect 417502 622658 417586 622894
rect 417822 622658 417854 622894
rect 417234 622574 417854 622658
rect 417234 622338 417266 622574
rect 417502 622338 417586 622574
rect 417822 622338 417854 622574
rect 417234 588894 417854 622338
rect 417234 588658 417266 588894
rect 417502 588658 417586 588894
rect 417822 588658 417854 588894
rect 417234 588574 417854 588658
rect 417234 588338 417266 588574
rect 417502 588338 417586 588574
rect 417822 588338 417854 588574
rect 417234 554894 417854 588338
rect 417234 554658 417266 554894
rect 417502 554658 417586 554894
rect 417822 554658 417854 554894
rect 417234 554574 417854 554658
rect 417234 554338 417266 554574
rect 417502 554338 417586 554574
rect 417822 554338 417854 554574
rect 417234 520894 417854 554338
rect 417234 520658 417266 520894
rect 417502 520658 417586 520894
rect 417822 520658 417854 520894
rect 417234 520574 417854 520658
rect 417234 520338 417266 520574
rect 417502 520338 417586 520574
rect 417822 520338 417854 520574
rect 417234 486894 417854 520338
rect 417234 486658 417266 486894
rect 417502 486658 417586 486894
rect 417822 486658 417854 486894
rect 417234 486574 417854 486658
rect 417234 486338 417266 486574
rect 417502 486338 417586 486574
rect 417822 486338 417854 486574
rect 417234 452894 417854 486338
rect 417234 452658 417266 452894
rect 417502 452658 417586 452894
rect 417822 452658 417854 452894
rect 417234 452574 417854 452658
rect 417234 452338 417266 452574
rect 417502 452338 417586 452574
rect 417822 452338 417854 452574
rect 417234 418894 417854 452338
rect 417234 418658 417266 418894
rect 417502 418658 417586 418894
rect 417822 418658 417854 418894
rect 417234 418574 417854 418658
rect 417234 418338 417266 418574
rect 417502 418338 417586 418574
rect 417822 418338 417854 418574
rect 417234 384894 417854 418338
rect 417234 384658 417266 384894
rect 417502 384658 417586 384894
rect 417822 384658 417854 384894
rect 417234 384574 417854 384658
rect 417234 384338 417266 384574
rect 417502 384338 417586 384574
rect 417822 384338 417854 384574
rect 417234 350894 417854 384338
rect 417234 350658 417266 350894
rect 417502 350658 417586 350894
rect 417822 350658 417854 350894
rect 417234 350574 417854 350658
rect 417234 350338 417266 350574
rect 417502 350338 417586 350574
rect 417822 350338 417854 350574
rect 417234 316894 417854 350338
rect 417234 316658 417266 316894
rect 417502 316658 417586 316894
rect 417822 316658 417854 316894
rect 417234 316574 417854 316658
rect 417234 316338 417266 316574
rect 417502 316338 417586 316574
rect 417822 316338 417854 316574
rect 417234 282894 417854 316338
rect 417234 282658 417266 282894
rect 417502 282658 417586 282894
rect 417822 282658 417854 282894
rect 417234 282574 417854 282658
rect 417234 282338 417266 282574
rect 417502 282338 417586 282574
rect 417822 282338 417854 282574
rect 417234 248894 417854 282338
rect 417234 248658 417266 248894
rect 417502 248658 417586 248894
rect 417822 248658 417854 248894
rect 417234 248574 417854 248658
rect 417234 248338 417266 248574
rect 417502 248338 417586 248574
rect 417822 248338 417854 248574
rect 417234 214894 417854 248338
rect 417234 214658 417266 214894
rect 417502 214658 417586 214894
rect 417822 214658 417854 214894
rect 417234 214574 417854 214658
rect 417234 214338 417266 214574
rect 417502 214338 417586 214574
rect 417822 214338 417854 214574
rect 417234 180894 417854 214338
rect 417234 180658 417266 180894
rect 417502 180658 417586 180894
rect 417822 180658 417854 180894
rect 417234 180574 417854 180658
rect 417234 180338 417266 180574
rect 417502 180338 417586 180574
rect 417822 180338 417854 180574
rect 417234 146894 417854 180338
rect 417234 146658 417266 146894
rect 417502 146658 417586 146894
rect 417822 146658 417854 146894
rect 417234 146574 417854 146658
rect 417234 146338 417266 146574
rect 417502 146338 417586 146574
rect 417822 146338 417854 146574
rect 417234 112894 417854 146338
rect 417234 112658 417266 112894
rect 417502 112658 417586 112894
rect 417822 112658 417854 112894
rect 417234 112574 417854 112658
rect 417234 112338 417266 112574
rect 417502 112338 417586 112574
rect 417822 112338 417854 112574
rect 417234 78894 417854 112338
rect 417234 78658 417266 78894
rect 417502 78658 417586 78894
rect 417822 78658 417854 78894
rect 417234 78574 417854 78658
rect 417234 78338 417266 78574
rect 417502 78338 417586 78574
rect 417822 78338 417854 78574
rect 417234 44894 417854 78338
rect 417234 44658 417266 44894
rect 417502 44658 417586 44894
rect 417822 44658 417854 44894
rect 417234 44574 417854 44658
rect 417234 44338 417266 44574
rect 417502 44338 417586 44574
rect 417822 44338 417854 44574
rect 417234 10894 417854 44338
rect 417234 10658 417266 10894
rect 417502 10658 417586 10894
rect 417822 10658 417854 10894
rect 417234 10574 417854 10658
rect 417234 10338 417266 10574
rect 417502 10338 417586 10574
rect 417822 10338 417854 10574
rect 417234 -2266 417854 10338
rect 417234 -2502 417266 -2266
rect 417502 -2502 417586 -2266
rect 417822 -2502 417854 -2266
rect 417234 -2586 417854 -2502
rect 417234 -2822 417266 -2586
rect 417502 -2822 417586 -2586
rect 417822 -2822 417854 -2586
rect 417234 -7654 417854 -2822
rect 420954 707718 421574 711590
rect 420954 707482 420986 707718
rect 421222 707482 421306 707718
rect 421542 707482 421574 707718
rect 420954 707398 421574 707482
rect 420954 707162 420986 707398
rect 421222 707162 421306 707398
rect 421542 707162 421574 707398
rect 420954 694614 421574 707162
rect 420954 694378 420986 694614
rect 421222 694378 421306 694614
rect 421542 694378 421574 694614
rect 420954 694294 421574 694378
rect 420954 694058 420986 694294
rect 421222 694058 421306 694294
rect 421542 694058 421574 694294
rect 420954 660614 421574 694058
rect 420954 660378 420986 660614
rect 421222 660378 421306 660614
rect 421542 660378 421574 660614
rect 420954 660294 421574 660378
rect 420954 660058 420986 660294
rect 421222 660058 421306 660294
rect 421542 660058 421574 660294
rect 420954 626614 421574 660058
rect 420954 626378 420986 626614
rect 421222 626378 421306 626614
rect 421542 626378 421574 626614
rect 420954 626294 421574 626378
rect 420954 626058 420986 626294
rect 421222 626058 421306 626294
rect 421542 626058 421574 626294
rect 420954 592614 421574 626058
rect 420954 592378 420986 592614
rect 421222 592378 421306 592614
rect 421542 592378 421574 592614
rect 420954 592294 421574 592378
rect 420954 592058 420986 592294
rect 421222 592058 421306 592294
rect 421542 592058 421574 592294
rect 420954 558614 421574 592058
rect 420954 558378 420986 558614
rect 421222 558378 421306 558614
rect 421542 558378 421574 558614
rect 420954 558294 421574 558378
rect 420954 558058 420986 558294
rect 421222 558058 421306 558294
rect 421542 558058 421574 558294
rect 420954 524614 421574 558058
rect 420954 524378 420986 524614
rect 421222 524378 421306 524614
rect 421542 524378 421574 524614
rect 420954 524294 421574 524378
rect 420954 524058 420986 524294
rect 421222 524058 421306 524294
rect 421542 524058 421574 524294
rect 420954 490614 421574 524058
rect 420954 490378 420986 490614
rect 421222 490378 421306 490614
rect 421542 490378 421574 490614
rect 420954 490294 421574 490378
rect 420954 490058 420986 490294
rect 421222 490058 421306 490294
rect 421542 490058 421574 490294
rect 420954 456614 421574 490058
rect 420954 456378 420986 456614
rect 421222 456378 421306 456614
rect 421542 456378 421574 456614
rect 420954 456294 421574 456378
rect 420954 456058 420986 456294
rect 421222 456058 421306 456294
rect 421542 456058 421574 456294
rect 420954 422614 421574 456058
rect 420954 422378 420986 422614
rect 421222 422378 421306 422614
rect 421542 422378 421574 422614
rect 420954 422294 421574 422378
rect 420954 422058 420986 422294
rect 421222 422058 421306 422294
rect 421542 422058 421574 422294
rect 420954 388614 421574 422058
rect 420954 388378 420986 388614
rect 421222 388378 421306 388614
rect 421542 388378 421574 388614
rect 420954 388294 421574 388378
rect 420954 388058 420986 388294
rect 421222 388058 421306 388294
rect 421542 388058 421574 388294
rect 420954 354614 421574 388058
rect 420954 354378 420986 354614
rect 421222 354378 421306 354614
rect 421542 354378 421574 354614
rect 420954 354294 421574 354378
rect 420954 354058 420986 354294
rect 421222 354058 421306 354294
rect 421542 354058 421574 354294
rect 420954 320614 421574 354058
rect 420954 320378 420986 320614
rect 421222 320378 421306 320614
rect 421542 320378 421574 320614
rect 420954 320294 421574 320378
rect 420954 320058 420986 320294
rect 421222 320058 421306 320294
rect 421542 320058 421574 320294
rect 420954 286614 421574 320058
rect 420954 286378 420986 286614
rect 421222 286378 421306 286614
rect 421542 286378 421574 286614
rect 420954 286294 421574 286378
rect 420954 286058 420986 286294
rect 421222 286058 421306 286294
rect 421542 286058 421574 286294
rect 420954 252614 421574 286058
rect 420954 252378 420986 252614
rect 421222 252378 421306 252614
rect 421542 252378 421574 252614
rect 420954 252294 421574 252378
rect 420954 252058 420986 252294
rect 421222 252058 421306 252294
rect 421542 252058 421574 252294
rect 420954 218614 421574 252058
rect 420954 218378 420986 218614
rect 421222 218378 421306 218614
rect 421542 218378 421574 218614
rect 420954 218294 421574 218378
rect 420954 218058 420986 218294
rect 421222 218058 421306 218294
rect 421542 218058 421574 218294
rect 420954 184614 421574 218058
rect 420954 184378 420986 184614
rect 421222 184378 421306 184614
rect 421542 184378 421574 184614
rect 420954 184294 421574 184378
rect 420954 184058 420986 184294
rect 421222 184058 421306 184294
rect 421542 184058 421574 184294
rect 420954 150614 421574 184058
rect 420954 150378 420986 150614
rect 421222 150378 421306 150614
rect 421542 150378 421574 150614
rect 420954 150294 421574 150378
rect 420954 150058 420986 150294
rect 421222 150058 421306 150294
rect 421542 150058 421574 150294
rect 420954 116614 421574 150058
rect 420954 116378 420986 116614
rect 421222 116378 421306 116614
rect 421542 116378 421574 116614
rect 420954 116294 421574 116378
rect 420954 116058 420986 116294
rect 421222 116058 421306 116294
rect 421542 116058 421574 116294
rect 420954 82614 421574 116058
rect 420954 82378 420986 82614
rect 421222 82378 421306 82614
rect 421542 82378 421574 82614
rect 420954 82294 421574 82378
rect 420954 82058 420986 82294
rect 421222 82058 421306 82294
rect 421542 82058 421574 82294
rect 420954 48614 421574 82058
rect 420954 48378 420986 48614
rect 421222 48378 421306 48614
rect 421542 48378 421574 48614
rect 420954 48294 421574 48378
rect 420954 48058 420986 48294
rect 421222 48058 421306 48294
rect 421542 48058 421574 48294
rect 420954 14614 421574 48058
rect 420954 14378 420986 14614
rect 421222 14378 421306 14614
rect 421542 14378 421574 14614
rect 420954 14294 421574 14378
rect 420954 14058 420986 14294
rect 421222 14058 421306 14294
rect 421542 14058 421574 14294
rect 420954 -3226 421574 14058
rect 420954 -3462 420986 -3226
rect 421222 -3462 421306 -3226
rect 421542 -3462 421574 -3226
rect 420954 -3546 421574 -3462
rect 420954 -3782 420986 -3546
rect 421222 -3782 421306 -3546
rect 421542 -3782 421574 -3546
rect 420954 -7654 421574 -3782
rect 424674 708678 425294 711590
rect 424674 708442 424706 708678
rect 424942 708442 425026 708678
rect 425262 708442 425294 708678
rect 424674 708358 425294 708442
rect 424674 708122 424706 708358
rect 424942 708122 425026 708358
rect 425262 708122 425294 708358
rect 424674 698334 425294 708122
rect 424674 698098 424706 698334
rect 424942 698098 425026 698334
rect 425262 698098 425294 698334
rect 424674 698014 425294 698098
rect 424674 697778 424706 698014
rect 424942 697778 425026 698014
rect 425262 697778 425294 698014
rect 424674 664334 425294 697778
rect 424674 664098 424706 664334
rect 424942 664098 425026 664334
rect 425262 664098 425294 664334
rect 424674 664014 425294 664098
rect 424674 663778 424706 664014
rect 424942 663778 425026 664014
rect 425262 663778 425294 664014
rect 424674 630334 425294 663778
rect 424674 630098 424706 630334
rect 424942 630098 425026 630334
rect 425262 630098 425294 630334
rect 424674 630014 425294 630098
rect 424674 629778 424706 630014
rect 424942 629778 425026 630014
rect 425262 629778 425294 630014
rect 424674 596334 425294 629778
rect 424674 596098 424706 596334
rect 424942 596098 425026 596334
rect 425262 596098 425294 596334
rect 424674 596014 425294 596098
rect 424674 595778 424706 596014
rect 424942 595778 425026 596014
rect 425262 595778 425294 596014
rect 424674 562334 425294 595778
rect 424674 562098 424706 562334
rect 424942 562098 425026 562334
rect 425262 562098 425294 562334
rect 424674 562014 425294 562098
rect 424674 561778 424706 562014
rect 424942 561778 425026 562014
rect 425262 561778 425294 562014
rect 424674 528334 425294 561778
rect 424674 528098 424706 528334
rect 424942 528098 425026 528334
rect 425262 528098 425294 528334
rect 424674 528014 425294 528098
rect 424674 527778 424706 528014
rect 424942 527778 425026 528014
rect 425262 527778 425294 528014
rect 424674 494334 425294 527778
rect 424674 494098 424706 494334
rect 424942 494098 425026 494334
rect 425262 494098 425294 494334
rect 424674 494014 425294 494098
rect 424674 493778 424706 494014
rect 424942 493778 425026 494014
rect 425262 493778 425294 494014
rect 424674 460334 425294 493778
rect 424674 460098 424706 460334
rect 424942 460098 425026 460334
rect 425262 460098 425294 460334
rect 424674 460014 425294 460098
rect 424674 459778 424706 460014
rect 424942 459778 425026 460014
rect 425262 459778 425294 460014
rect 424674 426334 425294 459778
rect 424674 426098 424706 426334
rect 424942 426098 425026 426334
rect 425262 426098 425294 426334
rect 424674 426014 425294 426098
rect 424674 425778 424706 426014
rect 424942 425778 425026 426014
rect 425262 425778 425294 426014
rect 424674 392334 425294 425778
rect 424674 392098 424706 392334
rect 424942 392098 425026 392334
rect 425262 392098 425294 392334
rect 424674 392014 425294 392098
rect 424674 391778 424706 392014
rect 424942 391778 425026 392014
rect 425262 391778 425294 392014
rect 424674 358334 425294 391778
rect 424674 358098 424706 358334
rect 424942 358098 425026 358334
rect 425262 358098 425294 358334
rect 424674 358014 425294 358098
rect 424674 357778 424706 358014
rect 424942 357778 425026 358014
rect 425262 357778 425294 358014
rect 424674 324334 425294 357778
rect 424674 324098 424706 324334
rect 424942 324098 425026 324334
rect 425262 324098 425294 324334
rect 424674 324014 425294 324098
rect 424674 323778 424706 324014
rect 424942 323778 425026 324014
rect 425262 323778 425294 324014
rect 424674 290334 425294 323778
rect 424674 290098 424706 290334
rect 424942 290098 425026 290334
rect 425262 290098 425294 290334
rect 424674 290014 425294 290098
rect 424674 289778 424706 290014
rect 424942 289778 425026 290014
rect 425262 289778 425294 290014
rect 424674 256334 425294 289778
rect 424674 256098 424706 256334
rect 424942 256098 425026 256334
rect 425262 256098 425294 256334
rect 424674 256014 425294 256098
rect 424674 255778 424706 256014
rect 424942 255778 425026 256014
rect 425262 255778 425294 256014
rect 424674 222334 425294 255778
rect 424674 222098 424706 222334
rect 424942 222098 425026 222334
rect 425262 222098 425294 222334
rect 424674 222014 425294 222098
rect 424674 221778 424706 222014
rect 424942 221778 425026 222014
rect 425262 221778 425294 222014
rect 424674 188334 425294 221778
rect 424674 188098 424706 188334
rect 424942 188098 425026 188334
rect 425262 188098 425294 188334
rect 424674 188014 425294 188098
rect 424674 187778 424706 188014
rect 424942 187778 425026 188014
rect 425262 187778 425294 188014
rect 424674 154334 425294 187778
rect 424674 154098 424706 154334
rect 424942 154098 425026 154334
rect 425262 154098 425294 154334
rect 424674 154014 425294 154098
rect 424674 153778 424706 154014
rect 424942 153778 425026 154014
rect 425262 153778 425294 154014
rect 424674 120334 425294 153778
rect 424674 120098 424706 120334
rect 424942 120098 425026 120334
rect 425262 120098 425294 120334
rect 424674 120014 425294 120098
rect 424674 119778 424706 120014
rect 424942 119778 425026 120014
rect 425262 119778 425294 120014
rect 424674 86334 425294 119778
rect 424674 86098 424706 86334
rect 424942 86098 425026 86334
rect 425262 86098 425294 86334
rect 424674 86014 425294 86098
rect 424674 85778 424706 86014
rect 424942 85778 425026 86014
rect 425262 85778 425294 86014
rect 424674 52334 425294 85778
rect 424674 52098 424706 52334
rect 424942 52098 425026 52334
rect 425262 52098 425294 52334
rect 424674 52014 425294 52098
rect 424674 51778 424706 52014
rect 424942 51778 425026 52014
rect 425262 51778 425294 52014
rect 424674 18334 425294 51778
rect 424674 18098 424706 18334
rect 424942 18098 425026 18334
rect 425262 18098 425294 18334
rect 424674 18014 425294 18098
rect 424674 17778 424706 18014
rect 424942 17778 425026 18014
rect 425262 17778 425294 18014
rect 424674 -4186 425294 17778
rect 424674 -4422 424706 -4186
rect 424942 -4422 425026 -4186
rect 425262 -4422 425294 -4186
rect 424674 -4506 425294 -4422
rect 424674 -4742 424706 -4506
rect 424942 -4742 425026 -4506
rect 425262 -4742 425294 -4506
rect 424674 -7654 425294 -4742
rect 428394 709638 429014 711590
rect 428394 709402 428426 709638
rect 428662 709402 428746 709638
rect 428982 709402 429014 709638
rect 428394 709318 429014 709402
rect 428394 709082 428426 709318
rect 428662 709082 428746 709318
rect 428982 709082 429014 709318
rect 428394 668054 429014 709082
rect 428394 667818 428426 668054
rect 428662 667818 428746 668054
rect 428982 667818 429014 668054
rect 428394 667734 429014 667818
rect 428394 667498 428426 667734
rect 428662 667498 428746 667734
rect 428982 667498 429014 667734
rect 428394 634054 429014 667498
rect 428394 633818 428426 634054
rect 428662 633818 428746 634054
rect 428982 633818 429014 634054
rect 428394 633734 429014 633818
rect 428394 633498 428426 633734
rect 428662 633498 428746 633734
rect 428982 633498 429014 633734
rect 428394 600054 429014 633498
rect 428394 599818 428426 600054
rect 428662 599818 428746 600054
rect 428982 599818 429014 600054
rect 428394 599734 429014 599818
rect 428394 599498 428426 599734
rect 428662 599498 428746 599734
rect 428982 599498 429014 599734
rect 428394 566054 429014 599498
rect 428394 565818 428426 566054
rect 428662 565818 428746 566054
rect 428982 565818 429014 566054
rect 428394 565734 429014 565818
rect 428394 565498 428426 565734
rect 428662 565498 428746 565734
rect 428982 565498 429014 565734
rect 428394 532054 429014 565498
rect 428394 531818 428426 532054
rect 428662 531818 428746 532054
rect 428982 531818 429014 532054
rect 428394 531734 429014 531818
rect 428394 531498 428426 531734
rect 428662 531498 428746 531734
rect 428982 531498 429014 531734
rect 428394 498054 429014 531498
rect 428394 497818 428426 498054
rect 428662 497818 428746 498054
rect 428982 497818 429014 498054
rect 428394 497734 429014 497818
rect 428394 497498 428426 497734
rect 428662 497498 428746 497734
rect 428982 497498 429014 497734
rect 428394 464054 429014 497498
rect 428394 463818 428426 464054
rect 428662 463818 428746 464054
rect 428982 463818 429014 464054
rect 428394 463734 429014 463818
rect 428394 463498 428426 463734
rect 428662 463498 428746 463734
rect 428982 463498 429014 463734
rect 428394 430054 429014 463498
rect 428394 429818 428426 430054
rect 428662 429818 428746 430054
rect 428982 429818 429014 430054
rect 428394 429734 429014 429818
rect 428394 429498 428426 429734
rect 428662 429498 428746 429734
rect 428982 429498 429014 429734
rect 428394 396054 429014 429498
rect 428394 395818 428426 396054
rect 428662 395818 428746 396054
rect 428982 395818 429014 396054
rect 428394 395734 429014 395818
rect 428394 395498 428426 395734
rect 428662 395498 428746 395734
rect 428982 395498 429014 395734
rect 428394 362054 429014 395498
rect 428394 361818 428426 362054
rect 428662 361818 428746 362054
rect 428982 361818 429014 362054
rect 428394 361734 429014 361818
rect 428394 361498 428426 361734
rect 428662 361498 428746 361734
rect 428982 361498 429014 361734
rect 428394 328054 429014 361498
rect 428394 327818 428426 328054
rect 428662 327818 428746 328054
rect 428982 327818 429014 328054
rect 428394 327734 429014 327818
rect 428394 327498 428426 327734
rect 428662 327498 428746 327734
rect 428982 327498 429014 327734
rect 428394 294054 429014 327498
rect 428394 293818 428426 294054
rect 428662 293818 428746 294054
rect 428982 293818 429014 294054
rect 428394 293734 429014 293818
rect 428394 293498 428426 293734
rect 428662 293498 428746 293734
rect 428982 293498 429014 293734
rect 428394 260054 429014 293498
rect 428394 259818 428426 260054
rect 428662 259818 428746 260054
rect 428982 259818 429014 260054
rect 428394 259734 429014 259818
rect 428394 259498 428426 259734
rect 428662 259498 428746 259734
rect 428982 259498 429014 259734
rect 428394 226054 429014 259498
rect 428394 225818 428426 226054
rect 428662 225818 428746 226054
rect 428982 225818 429014 226054
rect 428394 225734 429014 225818
rect 428394 225498 428426 225734
rect 428662 225498 428746 225734
rect 428982 225498 429014 225734
rect 428394 192054 429014 225498
rect 428394 191818 428426 192054
rect 428662 191818 428746 192054
rect 428982 191818 429014 192054
rect 428394 191734 429014 191818
rect 428394 191498 428426 191734
rect 428662 191498 428746 191734
rect 428982 191498 429014 191734
rect 428394 158054 429014 191498
rect 428394 157818 428426 158054
rect 428662 157818 428746 158054
rect 428982 157818 429014 158054
rect 428394 157734 429014 157818
rect 428394 157498 428426 157734
rect 428662 157498 428746 157734
rect 428982 157498 429014 157734
rect 428394 124054 429014 157498
rect 428394 123818 428426 124054
rect 428662 123818 428746 124054
rect 428982 123818 429014 124054
rect 428394 123734 429014 123818
rect 428394 123498 428426 123734
rect 428662 123498 428746 123734
rect 428982 123498 429014 123734
rect 428394 90054 429014 123498
rect 428394 89818 428426 90054
rect 428662 89818 428746 90054
rect 428982 89818 429014 90054
rect 428394 89734 429014 89818
rect 428394 89498 428426 89734
rect 428662 89498 428746 89734
rect 428982 89498 429014 89734
rect 428394 56054 429014 89498
rect 428394 55818 428426 56054
rect 428662 55818 428746 56054
rect 428982 55818 429014 56054
rect 428394 55734 429014 55818
rect 428394 55498 428426 55734
rect 428662 55498 428746 55734
rect 428982 55498 429014 55734
rect 428394 22054 429014 55498
rect 428394 21818 428426 22054
rect 428662 21818 428746 22054
rect 428982 21818 429014 22054
rect 428394 21734 429014 21818
rect 428394 21498 428426 21734
rect 428662 21498 428746 21734
rect 428982 21498 429014 21734
rect 428394 -5146 429014 21498
rect 428394 -5382 428426 -5146
rect 428662 -5382 428746 -5146
rect 428982 -5382 429014 -5146
rect 428394 -5466 429014 -5382
rect 428394 -5702 428426 -5466
rect 428662 -5702 428746 -5466
rect 428982 -5702 429014 -5466
rect 428394 -7654 429014 -5702
rect 432114 710598 432734 711590
rect 432114 710362 432146 710598
rect 432382 710362 432466 710598
rect 432702 710362 432734 710598
rect 432114 710278 432734 710362
rect 432114 710042 432146 710278
rect 432382 710042 432466 710278
rect 432702 710042 432734 710278
rect 432114 671774 432734 710042
rect 432114 671538 432146 671774
rect 432382 671538 432466 671774
rect 432702 671538 432734 671774
rect 432114 671454 432734 671538
rect 432114 671218 432146 671454
rect 432382 671218 432466 671454
rect 432702 671218 432734 671454
rect 432114 637774 432734 671218
rect 432114 637538 432146 637774
rect 432382 637538 432466 637774
rect 432702 637538 432734 637774
rect 432114 637454 432734 637538
rect 432114 637218 432146 637454
rect 432382 637218 432466 637454
rect 432702 637218 432734 637454
rect 432114 603774 432734 637218
rect 432114 603538 432146 603774
rect 432382 603538 432466 603774
rect 432702 603538 432734 603774
rect 432114 603454 432734 603538
rect 432114 603218 432146 603454
rect 432382 603218 432466 603454
rect 432702 603218 432734 603454
rect 432114 569774 432734 603218
rect 432114 569538 432146 569774
rect 432382 569538 432466 569774
rect 432702 569538 432734 569774
rect 432114 569454 432734 569538
rect 432114 569218 432146 569454
rect 432382 569218 432466 569454
rect 432702 569218 432734 569454
rect 432114 535774 432734 569218
rect 432114 535538 432146 535774
rect 432382 535538 432466 535774
rect 432702 535538 432734 535774
rect 432114 535454 432734 535538
rect 432114 535218 432146 535454
rect 432382 535218 432466 535454
rect 432702 535218 432734 535454
rect 432114 501774 432734 535218
rect 432114 501538 432146 501774
rect 432382 501538 432466 501774
rect 432702 501538 432734 501774
rect 432114 501454 432734 501538
rect 432114 501218 432146 501454
rect 432382 501218 432466 501454
rect 432702 501218 432734 501454
rect 432114 467774 432734 501218
rect 432114 467538 432146 467774
rect 432382 467538 432466 467774
rect 432702 467538 432734 467774
rect 432114 467454 432734 467538
rect 432114 467218 432146 467454
rect 432382 467218 432466 467454
rect 432702 467218 432734 467454
rect 432114 433774 432734 467218
rect 432114 433538 432146 433774
rect 432382 433538 432466 433774
rect 432702 433538 432734 433774
rect 432114 433454 432734 433538
rect 432114 433218 432146 433454
rect 432382 433218 432466 433454
rect 432702 433218 432734 433454
rect 432114 399774 432734 433218
rect 432114 399538 432146 399774
rect 432382 399538 432466 399774
rect 432702 399538 432734 399774
rect 432114 399454 432734 399538
rect 432114 399218 432146 399454
rect 432382 399218 432466 399454
rect 432702 399218 432734 399454
rect 432114 365774 432734 399218
rect 432114 365538 432146 365774
rect 432382 365538 432466 365774
rect 432702 365538 432734 365774
rect 432114 365454 432734 365538
rect 432114 365218 432146 365454
rect 432382 365218 432466 365454
rect 432702 365218 432734 365454
rect 432114 331774 432734 365218
rect 432114 331538 432146 331774
rect 432382 331538 432466 331774
rect 432702 331538 432734 331774
rect 432114 331454 432734 331538
rect 432114 331218 432146 331454
rect 432382 331218 432466 331454
rect 432702 331218 432734 331454
rect 432114 297774 432734 331218
rect 432114 297538 432146 297774
rect 432382 297538 432466 297774
rect 432702 297538 432734 297774
rect 432114 297454 432734 297538
rect 432114 297218 432146 297454
rect 432382 297218 432466 297454
rect 432702 297218 432734 297454
rect 432114 263774 432734 297218
rect 432114 263538 432146 263774
rect 432382 263538 432466 263774
rect 432702 263538 432734 263774
rect 432114 263454 432734 263538
rect 432114 263218 432146 263454
rect 432382 263218 432466 263454
rect 432702 263218 432734 263454
rect 432114 229774 432734 263218
rect 432114 229538 432146 229774
rect 432382 229538 432466 229774
rect 432702 229538 432734 229774
rect 432114 229454 432734 229538
rect 432114 229218 432146 229454
rect 432382 229218 432466 229454
rect 432702 229218 432734 229454
rect 432114 195774 432734 229218
rect 432114 195538 432146 195774
rect 432382 195538 432466 195774
rect 432702 195538 432734 195774
rect 432114 195454 432734 195538
rect 432114 195218 432146 195454
rect 432382 195218 432466 195454
rect 432702 195218 432734 195454
rect 432114 161774 432734 195218
rect 432114 161538 432146 161774
rect 432382 161538 432466 161774
rect 432702 161538 432734 161774
rect 432114 161454 432734 161538
rect 432114 161218 432146 161454
rect 432382 161218 432466 161454
rect 432702 161218 432734 161454
rect 432114 127774 432734 161218
rect 432114 127538 432146 127774
rect 432382 127538 432466 127774
rect 432702 127538 432734 127774
rect 432114 127454 432734 127538
rect 432114 127218 432146 127454
rect 432382 127218 432466 127454
rect 432702 127218 432734 127454
rect 432114 93774 432734 127218
rect 432114 93538 432146 93774
rect 432382 93538 432466 93774
rect 432702 93538 432734 93774
rect 432114 93454 432734 93538
rect 432114 93218 432146 93454
rect 432382 93218 432466 93454
rect 432702 93218 432734 93454
rect 432114 59774 432734 93218
rect 432114 59538 432146 59774
rect 432382 59538 432466 59774
rect 432702 59538 432734 59774
rect 432114 59454 432734 59538
rect 432114 59218 432146 59454
rect 432382 59218 432466 59454
rect 432702 59218 432734 59454
rect 432114 25774 432734 59218
rect 432114 25538 432146 25774
rect 432382 25538 432466 25774
rect 432702 25538 432734 25774
rect 432114 25454 432734 25538
rect 432114 25218 432146 25454
rect 432382 25218 432466 25454
rect 432702 25218 432734 25454
rect 432114 -6106 432734 25218
rect 432114 -6342 432146 -6106
rect 432382 -6342 432466 -6106
rect 432702 -6342 432734 -6106
rect 432114 -6426 432734 -6342
rect 432114 -6662 432146 -6426
rect 432382 -6662 432466 -6426
rect 432702 -6662 432734 -6426
rect 432114 -7654 432734 -6662
rect 435834 711558 436454 711590
rect 435834 711322 435866 711558
rect 436102 711322 436186 711558
rect 436422 711322 436454 711558
rect 435834 711238 436454 711322
rect 435834 711002 435866 711238
rect 436102 711002 436186 711238
rect 436422 711002 436454 711238
rect 435834 675494 436454 711002
rect 435834 675258 435866 675494
rect 436102 675258 436186 675494
rect 436422 675258 436454 675494
rect 435834 675174 436454 675258
rect 435834 674938 435866 675174
rect 436102 674938 436186 675174
rect 436422 674938 436454 675174
rect 435834 641494 436454 674938
rect 435834 641258 435866 641494
rect 436102 641258 436186 641494
rect 436422 641258 436454 641494
rect 435834 641174 436454 641258
rect 435834 640938 435866 641174
rect 436102 640938 436186 641174
rect 436422 640938 436454 641174
rect 435834 607494 436454 640938
rect 435834 607258 435866 607494
rect 436102 607258 436186 607494
rect 436422 607258 436454 607494
rect 435834 607174 436454 607258
rect 435834 606938 435866 607174
rect 436102 606938 436186 607174
rect 436422 606938 436454 607174
rect 435834 573494 436454 606938
rect 435834 573258 435866 573494
rect 436102 573258 436186 573494
rect 436422 573258 436454 573494
rect 435834 573174 436454 573258
rect 435834 572938 435866 573174
rect 436102 572938 436186 573174
rect 436422 572938 436454 573174
rect 435834 539494 436454 572938
rect 435834 539258 435866 539494
rect 436102 539258 436186 539494
rect 436422 539258 436454 539494
rect 435834 539174 436454 539258
rect 435834 538938 435866 539174
rect 436102 538938 436186 539174
rect 436422 538938 436454 539174
rect 435834 505494 436454 538938
rect 435834 505258 435866 505494
rect 436102 505258 436186 505494
rect 436422 505258 436454 505494
rect 435834 505174 436454 505258
rect 435834 504938 435866 505174
rect 436102 504938 436186 505174
rect 436422 504938 436454 505174
rect 435834 471494 436454 504938
rect 435834 471258 435866 471494
rect 436102 471258 436186 471494
rect 436422 471258 436454 471494
rect 435834 471174 436454 471258
rect 435834 470938 435866 471174
rect 436102 470938 436186 471174
rect 436422 470938 436454 471174
rect 435834 437494 436454 470938
rect 435834 437258 435866 437494
rect 436102 437258 436186 437494
rect 436422 437258 436454 437494
rect 435834 437174 436454 437258
rect 435834 436938 435866 437174
rect 436102 436938 436186 437174
rect 436422 436938 436454 437174
rect 435834 403494 436454 436938
rect 435834 403258 435866 403494
rect 436102 403258 436186 403494
rect 436422 403258 436454 403494
rect 435834 403174 436454 403258
rect 435834 402938 435866 403174
rect 436102 402938 436186 403174
rect 436422 402938 436454 403174
rect 435834 369494 436454 402938
rect 435834 369258 435866 369494
rect 436102 369258 436186 369494
rect 436422 369258 436454 369494
rect 435834 369174 436454 369258
rect 435834 368938 435866 369174
rect 436102 368938 436186 369174
rect 436422 368938 436454 369174
rect 435834 335494 436454 368938
rect 435834 335258 435866 335494
rect 436102 335258 436186 335494
rect 436422 335258 436454 335494
rect 435834 335174 436454 335258
rect 435834 334938 435866 335174
rect 436102 334938 436186 335174
rect 436422 334938 436454 335174
rect 435834 301494 436454 334938
rect 435834 301258 435866 301494
rect 436102 301258 436186 301494
rect 436422 301258 436454 301494
rect 435834 301174 436454 301258
rect 435834 300938 435866 301174
rect 436102 300938 436186 301174
rect 436422 300938 436454 301174
rect 435834 267494 436454 300938
rect 435834 267258 435866 267494
rect 436102 267258 436186 267494
rect 436422 267258 436454 267494
rect 435834 267174 436454 267258
rect 435834 266938 435866 267174
rect 436102 266938 436186 267174
rect 436422 266938 436454 267174
rect 435834 233494 436454 266938
rect 435834 233258 435866 233494
rect 436102 233258 436186 233494
rect 436422 233258 436454 233494
rect 435834 233174 436454 233258
rect 435834 232938 435866 233174
rect 436102 232938 436186 233174
rect 436422 232938 436454 233174
rect 435834 199494 436454 232938
rect 435834 199258 435866 199494
rect 436102 199258 436186 199494
rect 436422 199258 436454 199494
rect 435834 199174 436454 199258
rect 435834 198938 435866 199174
rect 436102 198938 436186 199174
rect 436422 198938 436454 199174
rect 435834 165494 436454 198938
rect 435834 165258 435866 165494
rect 436102 165258 436186 165494
rect 436422 165258 436454 165494
rect 435834 165174 436454 165258
rect 435834 164938 435866 165174
rect 436102 164938 436186 165174
rect 436422 164938 436454 165174
rect 435834 131494 436454 164938
rect 435834 131258 435866 131494
rect 436102 131258 436186 131494
rect 436422 131258 436454 131494
rect 435834 131174 436454 131258
rect 435834 130938 435866 131174
rect 436102 130938 436186 131174
rect 436422 130938 436454 131174
rect 435834 97494 436454 130938
rect 435834 97258 435866 97494
rect 436102 97258 436186 97494
rect 436422 97258 436454 97494
rect 435834 97174 436454 97258
rect 435834 96938 435866 97174
rect 436102 96938 436186 97174
rect 436422 96938 436454 97174
rect 435834 63494 436454 96938
rect 435834 63258 435866 63494
rect 436102 63258 436186 63494
rect 436422 63258 436454 63494
rect 435834 63174 436454 63258
rect 435834 62938 435866 63174
rect 436102 62938 436186 63174
rect 436422 62938 436454 63174
rect 435834 29494 436454 62938
rect 435834 29258 435866 29494
rect 436102 29258 436186 29494
rect 436422 29258 436454 29494
rect 435834 29174 436454 29258
rect 435834 28938 435866 29174
rect 436102 28938 436186 29174
rect 436422 28938 436454 29174
rect 435834 -7066 436454 28938
rect 435834 -7302 435866 -7066
rect 436102 -7302 436186 -7066
rect 436422 -7302 436454 -7066
rect 435834 -7386 436454 -7302
rect 435834 -7622 435866 -7386
rect 436102 -7622 436186 -7386
rect 436422 -7622 436454 -7386
rect 435834 -7654 436454 -7622
rect 443794 704838 444414 711590
rect 443794 704602 443826 704838
rect 444062 704602 444146 704838
rect 444382 704602 444414 704838
rect 443794 704518 444414 704602
rect 443794 704282 443826 704518
rect 444062 704282 444146 704518
rect 444382 704282 444414 704518
rect 443794 683454 444414 704282
rect 443794 683218 443826 683454
rect 444062 683218 444146 683454
rect 444382 683218 444414 683454
rect 443794 683134 444414 683218
rect 443794 682898 443826 683134
rect 444062 682898 444146 683134
rect 444382 682898 444414 683134
rect 443794 649454 444414 682898
rect 443794 649218 443826 649454
rect 444062 649218 444146 649454
rect 444382 649218 444414 649454
rect 443794 649134 444414 649218
rect 443794 648898 443826 649134
rect 444062 648898 444146 649134
rect 444382 648898 444414 649134
rect 443794 615454 444414 648898
rect 443794 615218 443826 615454
rect 444062 615218 444146 615454
rect 444382 615218 444414 615454
rect 443794 615134 444414 615218
rect 443794 614898 443826 615134
rect 444062 614898 444146 615134
rect 444382 614898 444414 615134
rect 443794 581454 444414 614898
rect 443794 581218 443826 581454
rect 444062 581218 444146 581454
rect 444382 581218 444414 581454
rect 443794 581134 444414 581218
rect 443794 580898 443826 581134
rect 444062 580898 444146 581134
rect 444382 580898 444414 581134
rect 443794 547454 444414 580898
rect 443794 547218 443826 547454
rect 444062 547218 444146 547454
rect 444382 547218 444414 547454
rect 443794 547134 444414 547218
rect 443794 546898 443826 547134
rect 444062 546898 444146 547134
rect 444382 546898 444414 547134
rect 443794 513454 444414 546898
rect 443794 513218 443826 513454
rect 444062 513218 444146 513454
rect 444382 513218 444414 513454
rect 443794 513134 444414 513218
rect 443794 512898 443826 513134
rect 444062 512898 444146 513134
rect 444382 512898 444414 513134
rect 443794 479454 444414 512898
rect 443794 479218 443826 479454
rect 444062 479218 444146 479454
rect 444382 479218 444414 479454
rect 443794 479134 444414 479218
rect 443794 478898 443826 479134
rect 444062 478898 444146 479134
rect 444382 478898 444414 479134
rect 443794 445454 444414 478898
rect 443794 445218 443826 445454
rect 444062 445218 444146 445454
rect 444382 445218 444414 445454
rect 443794 445134 444414 445218
rect 443794 444898 443826 445134
rect 444062 444898 444146 445134
rect 444382 444898 444414 445134
rect 443794 411454 444414 444898
rect 443794 411218 443826 411454
rect 444062 411218 444146 411454
rect 444382 411218 444414 411454
rect 443794 411134 444414 411218
rect 443794 410898 443826 411134
rect 444062 410898 444146 411134
rect 444382 410898 444414 411134
rect 443794 377454 444414 410898
rect 443794 377218 443826 377454
rect 444062 377218 444146 377454
rect 444382 377218 444414 377454
rect 443794 377134 444414 377218
rect 443794 376898 443826 377134
rect 444062 376898 444146 377134
rect 444382 376898 444414 377134
rect 443794 343454 444414 376898
rect 443794 343218 443826 343454
rect 444062 343218 444146 343454
rect 444382 343218 444414 343454
rect 443794 343134 444414 343218
rect 443794 342898 443826 343134
rect 444062 342898 444146 343134
rect 444382 342898 444414 343134
rect 443794 309454 444414 342898
rect 443794 309218 443826 309454
rect 444062 309218 444146 309454
rect 444382 309218 444414 309454
rect 443794 309134 444414 309218
rect 443794 308898 443826 309134
rect 444062 308898 444146 309134
rect 444382 308898 444414 309134
rect 443794 275454 444414 308898
rect 443794 275218 443826 275454
rect 444062 275218 444146 275454
rect 444382 275218 444414 275454
rect 443794 275134 444414 275218
rect 443794 274898 443826 275134
rect 444062 274898 444146 275134
rect 444382 274898 444414 275134
rect 443794 241454 444414 274898
rect 443794 241218 443826 241454
rect 444062 241218 444146 241454
rect 444382 241218 444414 241454
rect 443794 241134 444414 241218
rect 443794 240898 443826 241134
rect 444062 240898 444146 241134
rect 444382 240898 444414 241134
rect 443794 207454 444414 240898
rect 443794 207218 443826 207454
rect 444062 207218 444146 207454
rect 444382 207218 444414 207454
rect 443794 207134 444414 207218
rect 443794 206898 443826 207134
rect 444062 206898 444146 207134
rect 444382 206898 444414 207134
rect 443794 173454 444414 206898
rect 443794 173218 443826 173454
rect 444062 173218 444146 173454
rect 444382 173218 444414 173454
rect 443794 173134 444414 173218
rect 443794 172898 443826 173134
rect 444062 172898 444146 173134
rect 444382 172898 444414 173134
rect 443794 139454 444414 172898
rect 443794 139218 443826 139454
rect 444062 139218 444146 139454
rect 444382 139218 444414 139454
rect 443794 139134 444414 139218
rect 443794 138898 443826 139134
rect 444062 138898 444146 139134
rect 444382 138898 444414 139134
rect 443794 105454 444414 138898
rect 443794 105218 443826 105454
rect 444062 105218 444146 105454
rect 444382 105218 444414 105454
rect 443794 105134 444414 105218
rect 443794 104898 443826 105134
rect 444062 104898 444146 105134
rect 444382 104898 444414 105134
rect 443794 71454 444414 104898
rect 443794 71218 443826 71454
rect 444062 71218 444146 71454
rect 444382 71218 444414 71454
rect 443794 71134 444414 71218
rect 443794 70898 443826 71134
rect 444062 70898 444146 71134
rect 444382 70898 444414 71134
rect 443794 37454 444414 70898
rect 443794 37218 443826 37454
rect 444062 37218 444146 37454
rect 444382 37218 444414 37454
rect 443794 37134 444414 37218
rect 443794 36898 443826 37134
rect 444062 36898 444146 37134
rect 444382 36898 444414 37134
rect 443794 3454 444414 36898
rect 443794 3218 443826 3454
rect 444062 3218 444146 3454
rect 444382 3218 444414 3454
rect 443794 3134 444414 3218
rect 443794 2898 443826 3134
rect 444062 2898 444146 3134
rect 444382 2898 444414 3134
rect 443794 -346 444414 2898
rect 443794 -582 443826 -346
rect 444062 -582 444146 -346
rect 444382 -582 444414 -346
rect 443794 -666 444414 -582
rect 443794 -902 443826 -666
rect 444062 -902 444146 -666
rect 444382 -902 444414 -666
rect 443794 -7654 444414 -902
rect 447514 705798 448134 711590
rect 447514 705562 447546 705798
rect 447782 705562 447866 705798
rect 448102 705562 448134 705798
rect 447514 705478 448134 705562
rect 447514 705242 447546 705478
rect 447782 705242 447866 705478
rect 448102 705242 448134 705478
rect 447514 687174 448134 705242
rect 447514 686938 447546 687174
rect 447782 686938 447866 687174
rect 448102 686938 448134 687174
rect 447514 686854 448134 686938
rect 447514 686618 447546 686854
rect 447782 686618 447866 686854
rect 448102 686618 448134 686854
rect 447514 653174 448134 686618
rect 447514 652938 447546 653174
rect 447782 652938 447866 653174
rect 448102 652938 448134 653174
rect 447514 652854 448134 652938
rect 447514 652618 447546 652854
rect 447782 652618 447866 652854
rect 448102 652618 448134 652854
rect 447514 619174 448134 652618
rect 447514 618938 447546 619174
rect 447782 618938 447866 619174
rect 448102 618938 448134 619174
rect 447514 618854 448134 618938
rect 447514 618618 447546 618854
rect 447782 618618 447866 618854
rect 448102 618618 448134 618854
rect 447514 585174 448134 618618
rect 447514 584938 447546 585174
rect 447782 584938 447866 585174
rect 448102 584938 448134 585174
rect 447514 584854 448134 584938
rect 447514 584618 447546 584854
rect 447782 584618 447866 584854
rect 448102 584618 448134 584854
rect 447514 551174 448134 584618
rect 447514 550938 447546 551174
rect 447782 550938 447866 551174
rect 448102 550938 448134 551174
rect 447514 550854 448134 550938
rect 447514 550618 447546 550854
rect 447782 550618 447866 550854
rect 448102 550618 448134 550854
rect 447514 517174 448134 550618
rect 447514 516938 447546 517174
rect 447782 516938 447866 517174
rect 448102 516938 448134 517174
rect 447514 516854 448134 516938
rect 447514 516618 447546 516854
rect 447782 516618 447866 516854
rect 448102 516618 448134 516854
rect 447514 483174 448134 516618
rect 447514 482938 447546 483174
rect 447782 482938 447866 483174
rect 448102 482938 448134 483174
rect 447514 482854 448134 482938
rect 447514 482618 447546 482854
rect 447782 482618 447866 482854
rect 448102 482618 448134 482854
rect 447514 449174 448134 482618
rect 447514 448938 447546 449174
rect 447782 448938 447866 449174
rect 448102 448938 448134 449174
rect 447514 448854 448134 448938
rect 447514 448618 447546 448854
rect 447782 448618 447866 448854
rect 448102 448618 448134 448854
rect 447514 415174 448134 448618
rect 447514 414938 447546 415174
rect 447782 414938 447866 415174
rect 448102 414938 448134 415174
rect 447514 414854 448134 414938
rect 447514 414618 447546 414854
rect 447782 414618 447866 414854
rect 448102 414618 448134 414854
rect 447514 381174 448134 414618
rect 447514 380938 447546 381174
rect 447782 380938 447866 381174
rect 448102 380938 448134 381174
rect 447514 380854 448134 380938
rect 447514 380618 447546 380854
rect 447782 380618 447866 380854
rect 448102 380618 448134 380854
rect 447514 347174 448134 380618
rect 447514 346938 447546 347174
rect 447782 346938 447866 347174
rect 448102 346938 448134 347174
rect 447514 346854 448134 346938
rect 447514 346618 447546 346854
rect 447782 346618 447866 346854
rect 448102 346618 448134 346854
rect 447514 313174 448134 346618
rect 447514 312938 447546 313174
rect 447782 312938 447866 313174
rect 448102 312938 448134 313174
rect 447514 312854 448134 312938
rect 447514 312618 447546 312854
rect 447782 312618 447866 312854
rect 448102 312618 448134 312854
rect 447514 279174 448134 312618
rect 447514 278938 447546 279174
rect 447782 278938 447866 279174
rect 448102 278938 448134 279174
rect 447514 278854 448134 278938
rect 447514 278618 447546 278854
rect 447782 278618 447866 278854
rect 448102 278618 448134 278854
rect 447514 245174 448134 278618
rect 447514 244938 447546 245174
rect 447782 244938 447866 245174
rect 448102 244938 448134 245174
rect 447514 244854 448134 244938
rect 447514 244618 447546 244854
rect 447782 244618 447866 244854
rect 448102 244618 448134 244854
rect 447514 211174 448134 244618
rect 447514 210938 447546 211174
rect 447782 210938 447866 211174
rect 448102 210938 448134 211174
rect 447514 210854 448134 210938
rect 447514 210618 447546 210854
rect 447782 210618 447866 210854
rect 448102 210618 448134 210854
rect 447514 177174 448134 210618
rect 447514 176938 447546 177174
rect 447782 176938 447866 177174
rect 448102 176938 448134 177174
rect 447514 176854 448134 176938
rect 447514 176618 447546 176854
rect 447782 176618 447866 176854
rect 448102 176618 448134 176854
rect 447514 143174 448134 176618
rect 447514 142938 447546 143174
rect 447782 142938 447866 143174
rect 448102 142938 448134 143174
rect 447514 142854 448134 142938
rect 447514 142618 447546 142854
rect 447782 142618 447866 142854
rect 448102 142618 448134 142854
rect 447514 109174 448134 142618
rect 447514 108938 447546 109174
rect 447782 108938 447866 109174
rect 448102 108938 448134 109174
rect 447514 108854 448134 108938
rect 447514 108618 447546 108854
rect 447782 108618 447866 108854
rect 448102 108618 448134 108854
rect 447514 75174 448134 108618
rect 447514 74938 447546 75174
rect 447782 74938 447866 75174
rect 448102 74938 448134 75174
rect 447514 74854 448134 74938
rect 447514 74618 447546 74854
rect 447782 74618 447866 74854
rect 448102 74618 448134 74854
rect 447514 41174 448134 74618
rect 447514 40938 447546 41174
rect 447782 40938 447866 41174
rect 448102 40938 448134 41174
rect 447514 40854 448134 40938
rect 447514 40618 447546 40854
rect 447782 40618 447866 40854
rect 448102 40618 448134 40854
rect 447514 7174 448134 40618
rect 447514 6938 447546 7174
rect 447782 6938 447866 7174
rect 448102 6938 448134 7174
rect 447514 6854 448134 6938
rect 447514 6618 447546 6854
rect 447782 6618 447866 6854
rect 448102 6618 448134 6854
rect 447514 -1306 448134 6618
rect 447514 -1542 447546 -1306
rect 447782 -1542 447866 -1306
rect 448102 -1542 448134 -1306
rect 447514 -1626 448134 -1542
rect 447514 -1862 447546 -1626
rect 447782 -1862 447866 -1626
rect 448102 -1862 448134 -1626
rect 447514 -7654 448134 -1862
rect 451234 706758 451854 711590
rect 451234 706522 451266 706758
rect 451502 706522 451586 706758
rect 451822 706522 451854 706758
rect 451234 706438 451854 706522
rect 451234 706202 451266 706438
rect 451502 706202 451586 706438
rect 451822 706202 451854 706438
rect 451234 690894 451854 706202
rect 451234 690658 451266 690894
rect 451502 690658 451586 690894
rect 451822 690658 451854 690894
rect 451234 690574 451854 690658
rect 451234 690338 451266 690574
rect 451502 690338 451586 690574
rect 451822 690338 451854 690574
rect 451234 656894 451854 690338
rect 451234 656658 451266 656894
rect 451502 656658 451586 656894
rect 451822 656658 451854 656894
rect 451234 656574 451854 656658
rect 451234 656338 451266 656574
rect 451502 656338 451586 656574
rect 451822 656338 451854 656574
rect 451234 622894 451854 656338
rect 451234 622658 451266 622894
rect 451502 622658 451586 622894
rect 451822 622658 451854 622894
rect 451234 622574 451854 622658
rect 451234 622338 451266 622574
rect 451502 622338 451586 622574
rect 451822 622338 451854 622574
rect 451234 588894 451854 622338
rect 451234 588658 451266 588894
rect 451502 588658 451586 588894
rect 451822 588658 451854 588894
rect 451234 588574 451854 588658
rect 451234 588338 451266 588574
rect 451502 588338 451586 588574
rect 451822 588338 451854 588574
rect 451234 554894 451854 588338
rect 451234 554658 451266 554894
rect 451502 554658 451586 554894
rect 451822 554658 451854 554894
rect 451234 554574 451854 554658
rect 451234 554338 451266 554574
rect 451502 554338 451586 554574
rect 451822 554338 451854 554574
rect 451234 520894 451854 554338
rect 451234 520658 451266 520894
rect 451502 520658 451586 520894
rect 451822 520658 451854 520894
rect 451234 520574 451854 520658
rect 451234 520338 451266 520574
rect 451502 520338 451586 520574
rect 451822 520338 451854 520574
rect 451234 486894 451854 520338
rect 451234 486658 451266 486894
rect 451502 486658 451586 486894
rect 451822 486658 451854 486894
rect 451234 486574 451854 486658
rect 451234 486338 451266 486574
rect 451502 486338 451586 486574
rect 451822 486338 451854 486574
rect 451234 452894 451854 486338
rect 451234 452658 451266 452894
rect 451502 452658 451586 452894
rect 451822 452658 451854 452894
rect 451234 452574 451854 452658
rect 451234 452338 451266 452574
rect 451502 452338 451586 452574
rect 451822 452338 451854 452574
rect 451234 418894 451854 452338
rect 451234 418658 451266 418894
rect 451502 418658 451586 418894
rect 451822 418658 451854 418894
rect 451234 418574 451854 418658
rect 451234 418338 451266 418574
rect 451502 418338 451586 418574
rect 451822 418338 451854 418574
rect 451234 384894 451854 418338
rect 451234 384658 451266 384894
rect 451502 384658 451586 384894
rect 451822 384658 451854 384894
rect 451234 384574 451854 384658
rect 451234 384338 451266 384574
rect 451502 384338 451586 384574
rect 451822 384338 451854 384574
rect 451234 350894 451854 384338
rect 451234 350658 451266 350894
rect 451502 350658 451586 350894
rect 451822 350658 451854 350894
rect 451234 350574 451854 350658
rect 451234 350338 451266 350574
rect 451502 350338 451586 350574
rect 451822 350338 451854 350574
rect 451234 316894 451854 350338
rect 451234 316658 451266 316894
rect 451502 316658 451586 316894
rect 451822 316658 451854 316894
rect 451234 316574 451854 316658
rect 451234 316338 451266 316574
rect 451502 316338 451586 316574
rect 451822 316338 451854 316574
rect 451234 282894 451854 316338
rect 451234 282658 451266 282894
rect 451502 282658 451586 282894
rect 451822 282658 451854 282894
rect 451234 282574 451854 282658
rect 451234 282338 451266 282574
rect 451502 282338 451586 282574
rect 451822 282338 451854 282574
rect 451234 248894 451854 282338
rect 451234 248658 451266 248894
rect 451502 248658 451586 248894
rect 451822 248658 451854 248894
rect 451234 248574 451854 248658
rect 451234 248338 451266 248574
rect 451502 248338 451586 248574
rect 451822 248338 451854 248574
rect 451234 214894 451854 248338
rect 451234 214658 451266 214894
rect 451502 214658 451586 214894
rect 451822 214658 451854 214894
rect 451234 214574 451854 214658
rect 451234 214338 451266 214574
rect 451502 214338 451586 214574
rect 451822 214338 451854 214574
rect 451234 180894 451854 214338
rect 451234 180658 451266 180894
rect 451502 180658 451586 180894
rect 451822 180658 451854 180894
rect 451234 180574 451854 180658
rect 451234 180338 451266 180574
rect 451502 180338 451586 180574
rect 451822 180338 451854 180574
rect 451234 146894 451854 180338
rect 451234 146658 451266 146894
rect 451502 146658 451586 146894
rect 451822 146658 451854 146894
rect 451234 146574 451854 146658
rect 451234 146338 451266 146574
rect 451502 146338 451586 146574
rect 451822 146338 451854 146574
rect 451234 112894 451854 146338
rect 451234 112658 451266 112894
rect 451502 112658 451586 112894
rect 451822 112658 451854 112894
rect 451234 112574 451854 112658
rect 451234 112338 451266 112574
rect 451502 112338 451586 112574
rect 451822 112338 451854 112574
rect 451234 78894 451854 112338
rect 451234 78658 451266 78894
rect 451502 78658 451586 78894
rect 451822 78658 451854 78894
rect 451234 78574 451854 78658
rect 451234 78338 451266 78574
rect 451502 78338 451586 78574
rect 451822 78338 451854 78574
rect 451234 44894 451854 78338
rect 451234 44658 451266 44894
rect 451502 44658 451586 44894
rect 451822 44658 451854 44894
rect 451234 44574 451854 44658
rect 451234 44338 451266 44574
rect 451502 44338 451586 44574
rect 451822 44338 451854 44574
rect 451234 10894 451854 44338
rect 451234 10658 451266 10894
rect 451502 10658 451586 10894
rect 451822 10658 451854 10894
rect 451234 10574 451854 10658
rect 451234 10338 451266 10574
rect 451502 10338 451586 10574
rect 451822 10338 451854 10574
rect 451234 -2266 451854 10338
rect 451234 -2502 451266 -2266
rect 451502 -2502 451586 -2266
rect 451822 -2502 451854 -2266
rect 451234 -2586 451854 -2502
rect 451234 -2822 451266 -2586
rect 451502 -2822 451586 -2586
rect 451822 -2822 451854 -2586
rect 451234 -7654 451854 -2822
rect 454954 707718 455574 711590
rect 454954 707482 454986 707718
rect 455222 707482 455306 707718
rect 455542 707482 455574 707718
rect 454954 707398 455574 707482
rect 454954 707162 454986 707398
rect 455222 707162 455306 707398
rect 455542 707162 455574 707398
rect 454954 694614 455574 707162
rect 454954 694378 454986 694614
rect 455222 694378 455306 694614
rect 455542 694378 455574 694614
rect 454954 694294 455574 694378
rect 454954 694058 454986 694294
rect 455222 694058 455306 694294
rect 455542 694058 455574 694294
rect 454954 660614 455574 694058
rect 454954 660378 454986 660614
rect 455222 660378 455306 660614
rect 455542 660378 455574 660614
rect 454954 660294 455574 660378
rect 454954 660058 454986 660294
rect 455222 660058 455306 660294
rect 455542 660058 455574 660294
rect 454954 626614 455574 660058
rect 454954 626378 454986 626614
rect 455222 626378 455306 626614
rect 455542 626378 455574 626614
rect 454954 626294 455574 626378
rect 454954 626058 454986 626294
rect 455222 626058 455306 626294
rect 455542 626058 455574 626294
rect 454954 592614 455574 626058
rect 454954 592378 454986 592614
rect 455222 592378 455306 592614
rect 455542 592378 455574 592614
rect 454954 592294 455574 592378
rect 454954 592058 454986 592294
rect 455222 592058 455306 592294
rect 455542 592058 455574 592294
rect 454954 558614 455574 592058
rect 454954 558378 454986 558614
rect 455222 558378 455306 558614
rect 455542 558378 455574 558614
rect 454954 558294 455574 558378
rect 454954 558058 454986 558294
rect 455222 558058 455306 558294
rect 455542 558058 455574 558294
rect 454954 524614 455574 558058
rect 454954 524378 454986 524614
rect 455222 524378 455306 524614
rect 455542 524378 455574 524614
rect 454954 524294 455574 524378
rect 454954 524058 454986 524294
rect 455222 524058 455306 524294
rect 455542 524058 455574 524294
rect 454954 490614 455574 524058
rect 454954 490378 454986 490614
rect 455222 490378 455306 490614
rect 455542 490378 455574 490614
rect 454954 490294 455574 490378
rect 454954 490058 454986 490294
rect 455222 490058 455306 490294
rect 455542 490058 455574 490294
rect 454954 456614 455574 490058
rect 454954 456378 454986 456614
rect 455222 456378 455306 456614
rect 455542 456378 455574 456614
rect 454954 456294 455574 456378
rect 454954 456058 454986 456294
rect 455222 456058 455306 456294
rect 455542 456058 455574 456294
rect 454954 422614 455574 456058
rect 454954 422378 454986 422614
rect 455222 422378 455306 422614
rect 455542 422378 455574 422614
rect 454954 422294 455574 422378
rect 454954 422058 454986 422294
rect 455222 422058 455306 422294
rect 455542 422058 455574 422294
rect 454954 388614 455574 422058
rect 454954 388378 454986 388614
rect 455222 388378 455306 388614
rect 455542 388378 455574 388614
rect 454954 388294 455574 388378
rect 454954 388058 454986 388294
rect 455222 388058 455306 388294
rect 455542 388058 455574 388294
rect 454954 354614 455574 388058
rect 454954 354378 454986 354614
rect 455222 354378 455306 354614
rect 455542 354378 455574 354614
rect 454954 354294 455574 354378
rect 454954 354058 454986 354294
rect 455222 354058 455306 354294
rect 455542 354058 455574 354294
rect 454954 320614 455574 354058
rect 454954 320378 454986 320614
rect 455222 320378 455306 320614
rect 455542 320378 455574 320614
rect 454954 320294 455574 320378
rect 454954 320058 454986 320294
rect 455222 320058 455306 320294
rect 455542 320058 455574 320294
rect 454954 286614 455574 320058
rect 454954 286378 454986 286614
rect 455222 286378 455306 286614
rect 455542 286378 455574 286614
rect 454954 286294 455574 286378
rect 454954 286058 454986 286294
rect 455222 286058 455306 286294
rect 455542 286058 455574 286294
rect 454954 252614 455574 286058
rect 454954 252378 454986 252614
rect 455222 252378 455306 252614
rect 455542 252378 455574 252614
rect 454954 252294 455574 252378
rect 454954 252058 454986 252294
rect 455222 252058 455306 252294
rect 455542 252058 455574 252294
rect 454954 218614 455574 252058
rect 454954 218378 454986 218614
rect 455222 218378 455306 218614
rect 455542 218378 455574 218614
rect 454954 218294 455574 218378
rect 454954 218058 454986 218294
rect 455222 218058 455306 218294
rect 455542 218058 455574 218294
rect 454954 184614 455574 218058
rect 454954 184378 454986 184614
rect 455222 184378 455306 184614
rect 455542 184378 455574 184614
rect 454954 184294 455574 184378
rect 454954 184058 454986 184294
rect 455222 184058 455306 184294
rect 455542 184058 455574 184294
rect 454954 150614 455574 184058
rect 454954 150378 454986 150614
rect 455222 150378 455306 150614
rect 455542 150378 455574 150614
rect 454954 150294 455574 150378
rect 454954 150058 454986 150294
rect 455222 150058 455306 150294
rect 455542 150058 455574 150294
rect 454954 116614 455574 150058
rect 454954 116378 454986 116614
rect 455222 116378 455306 116614
rect 455542 116378 455574 116614
rect 454954 116294 455574 116378
rect 454954 116058 454986 116294
rect 455222 116058 455306 116294
rect 455542 116058 455574 116294
rect 454954 82614 455574 116058
rect 454954 82378 454986 82614
rect 455222 82378 455306 82614
rect 455542 82378 455574 82614
rect 454954 82294 455574 82378
rect 454954 82058 454986 82294
rect 455222 82058 455306 82294
rect 455542 82058 455574 82294
rect 454954 48614 455574 82058
rect 454954 48378 454986 48614
rect 455222 48378 455306 48614
rect 455542 48378 455574 48614
rect 454954 48294 455574 48378
rect 454954 48058 454986 48294
rect 455222 48058 455306 48294
rect 455542 48058 455574 48294
rect 454954 14614 455574 48058
rect 454954 14378 454986 14614
rect 455222 14378 455306 14614
rect 455542 14378 455574 14614
rect 454954 14294 455574 14378
rect 454954 14058 454986 14294
rect 455222 14058 455306 14294
rect 455542 14058 455574 14294
rect 454954 -3226 455574 14058
rect 454954 -3462 454986 -3226
rect 455222 -3462 455306 -3226
rect 455542 -3462 455574 -3226
rect 454954 -3546 455574 -3462
rect 454954 -3782 454986 -3546
rect 455222 -3782 455306 -3546
rect 455542 -3782 455574 -3546
rect 454954 -7654 455574 -3782
rect 458674 708678 459294 711590
rect 458674 708442 458706 708678
rect 458942 708442 459026 708678
rect 459262 708442 459294 708678
rect 458674 708358 459294 708442
rect 458674 708122 458706 708358
rect 458942 708122 459026 708358
rect 459262 708122 459294 708358
rect 458674 698334 459294 708122
rect 458674 698098 458706 698334
rect 458942 698098 459026 698334
rect 459262 698098 459294 698334
rect 458674 698014 459294 698098
rect 458674 697778 458706 698014
rect 458942 697778 459026 698014
rect 459262 697778 459294 698014
rect 458674 664334 459294 697778
rect 458674 664098 458706 664334
rect 458942 664098 459026 664334
rect 459262 664098 459294 664334
rect 458674 664014 459294 664098
rect 458674 663778 458706 664014
rect 458942 663778 459026 664014
rect 459262 663778 459294 664014
rect 458674 630334 459294 663778
rect 458674 630098 458706 630334
rect 458942 630098 459026 630334
rect 459262 630098 459294 630334
rect 458674 630014 459294 630098
rect 458674 629778 458706 630014
rect 458942 629778 459026 630014
rect 459262 629778 459294 630014
rect 458674 596334 459294 629778
rect 458674 596098 458706 596334
rect 458942 596098 459026 596334
rect 459262 596098 459294 596334
rect 458674 596014 459294 596098
rect 458674 595778 458706 596014
rect 458942 595778 459026 596014
rect 459262 595778 459294 596014
rect 458674 562334 459294 595778
rect 458674 562098 458706 562334
rect 458942 562098 459026 562334
rect 459262 562098 459294 562334
rect 458674 562014 459294 562098
rect 458674 561778 458706 562014
rect 458942 561778 459026 562014
rect 459262 561778 459294 562014
rect 458674 528334 459294 561778
rect 458674 528098 458706 528334
rect 458942 528098 459026 528334
rect 459262 528098 459294 528334
rect 458674 528014 459294 528098
rect 458674 527778 458706 528014
rect 458942 527778 459026 528014
rect 459262 527778 459294 528014
rect 458674 494334 459294 527778
rect 458674 494098 458706 494334
rect 458942 494098 459026 494334
rect 459262 494098 459294 494334
rect 458674 494014 459294 494098
rect 458674 493778 458706 494014
rect 458942 493778 459026 494014
rect 459262 493778 459294 494014
rect 458674 460334 459294 493778
rect 458674 460098 458706 460334
rect 458942 460098 459026 460334
rect 459262 460098 459294 460334
rect 458674 460014 459294 460098
rect 458674 459778 458706 460014
rect 458942 459778 459026 460014
rect 459262 459778 459294 460014
rect 458674 426334 459294 459778
rect 458674 426098 458706 426334
rect 458942 426098 459026 426334
rect 459262 426098 459294 426334
rect 458674 426014 459294 426098
rect 458674 425778 458706 426014
rect 458942 425778 459026 426014
rect 459262 425778 459294 426014
rect 458674 392334 459294 425778
rect 458674 392098 458706 392334
rect 458942 392098 459026 392334
rect 459262 392098 459294 392334
rect 458674 392014 459294 392098
rect 458674 391778 458706 392014
rect 458942 391778 459026 392014
rect 459262 391778 459294 392014
rect 458674 358334 459294 391778
rect 458674 358098 458706 358334
rect 458942 358098 459026 358334
rect 459262 358098 459294 358334
rect 458674 358014 459294 358098
rect 458674 357778 458706 358014
rect 458942 357778 459026 358014
rect 459262 357778 459294 358014
rect 458674 324334 459294 357778
rect 458674 324098 458706 324334
rect 458942 324098 459026 324334
rect 459262 324098 459294 324334
rect 458674 324014 459294 324098
rect 458674 323778 458706 324014
rect 458942 323778 459026 324014
rect 459262 323778 459294 324014
rect 458674 290334 459294 323778
rect 458674 290098 458706 290334
rect 458942 290098 459026 290334
rect 459262 290098 459294 290334
rect 458674 290014 459294 290098
rect 458674 289778 458706 290014
rect 458942 289778 459026 290014
rect 459262 289778 459294 290014
rect 458674 256334 459294 289778
rect 458674 256098 458706 256334
rect 458942 256098 459026 256334
rect 459262 256098 459294 256334
rect 458674 256014 459294 256098
rect 458674 255778 458706 256014
rect 458942 255778 459026 256014
rect 459262 255778 459294 256014
rect 458674 222334 459294 255778
rect 458674 222098 458706 222334
rect 458942 222098 459026 222334
rect 459262 222098 459294 222334
rect 458674 222014 459294 222098
rect 458674 221778 458706 222014
rect 458942 221778 459026 222014
rect 459262 221778 459294 222014
rect 458674 188334 459294 221778
rect 458674 188098 458706 188334
rect 458942 188098 459026 188334
rect 459262 188098 459294 188334
rect 458674 188014 459294 188098
rect 458674 187778 458706 188014
rect 458942 187778 459026 188014
rect 459262 187778 459294 188014
rect 458674 154334 459294 187778
rect 458674 154098 458706 154334
rect 458942 154098 459026 154334
rect 459262 154098 459294 154334
rect 458674 154014 459294 154098
rect 458674 153778 458706 154014
rect 458942 153778 459026 154014
rect 459262 153778 459294 154014
rect 458674 120334 459294 153778
rect 458674 120098 458706 120334
rect 458942 120098 459026 120334
rect 459262 120098 459294 120334
rect 458674 120014 459294 120098
rect 458674 119778 458706 120014
rect 458942 119778 459026 120014
rect 459262 119778 459294 120014
rect 458674 86334 459294 119778
rect 458674 86098 458706 86334
rect 458942 86098 459026 86334
rect 459262 86098 459294 86334
rect 458674 86014 459294 86098
rect 458674 85778 458706 86014
rect 458942 85778 459026 86014
rect 459262 85778 459294 86014
rect 458674 52334 459294 85778
rect 458674 52098 458706 52334
rect 458942 52098 459026 52334
rect 459262 52098 459294 52334
rect 458674 52014 459294 52098
rect 458674 51778 458706 52014
rect 458942 51778 459026 52014
rect 459262 51778 459294 52014
rect 458674 18334 459294 51778
rect 458674 18098 458706 18334
rect 458942 18098 459026 18334
rect 459262 18098 459294 18334
rect 458674 18014 459294 18098
rect 458674 17778 458706 18014
rect 458942 17778 459026 18014
rect 459262 17778 459294 18014
rect 458674 -4186 459294 17778
rect 458674 -4422 458706 -4186
rect 458942 -4422 459026 -4186
rect 459262 -4422 459294 -4186
rect 458674 -4506 459294 -4422
rect 458674 -4742 458706 -4506
rect 458942 -4742 459026 -4506
rect 459262 -4742 459294 -4506
rect 458674 -7654 459294 -4742
rect 462394 709638 463014 711590
rect 462394 709402 462426 709638
rect 462662 709402 462746 709638
rect 462982 709402 463014 709638
rect 462394 709318 463014 709402
rect 462394 709082 462426 709318
rect 462662 709082 462746 709318
rect 462982 709082 463014 709318
rect 462394 668054 463014 709082
rect 462394 667818 462426 668054
rect 462662 667818 462746 668054
rect 462982 667818 463014 668054
rect 462394 667734 463014 667818
rect 462394 667498 462426 667734
rect 462662 667498 462746 667734
rect 462982 667498 463014 667734
rect 462394 634054 463014 667498
rect 462394 633818 462426 634054
rect 462662 633818 462746 634054
rect 462982 633818 463014 634054
rect 462394 633734 463014 633818
rect 462394 633498 462426 633734
rect 462662 633498 462746 633734
rect 462982 633498 463014 633734
rect 462394 600054 463014 633498
rect 462394 599818 462426 600054
rect 462662 599818 462746 600054
rect 462982 599818 463014 600054
rect 462394 599734 463014 599818
rect 462394 599498 462426 599734
rect 462662 599498 462746 599734
rect 462982 599498 463014 599734
rect 462394 566054 463014 599498
rect 462394 565818 462426 566054
rect 462662 565818 462746 566054
rect 462982 565818 463014 566054
rect 462394 565734 463014 565818
rect 462394 565498 462426 565734
rect 462662 565498 462746 565734
rect 462982 565498 463014 565734
rect 462394 532054 463014 565498
rect 462394 531818 462426 532054
rect 462662 531818 462746 532054
rect 462982 531818 463014 532054
rect 462394 531734 463014 531818
rect 462394 531498 462426 531734
rect 462662 531498 462746 531734
rect 462982 531498 463014 531734
rect 462394 498054 463014 531498
rect 462394 497818 462426 498054
rect 462662 497818 462746 498054
rect 462982 497818 463014 498054
rect 462394 497734 463014 497818
rect 462394 497498 462426 497734
rect 462662 497498 462746 497734
rect 462982 497498 463014 497734
rect 462394 464054 463014 497498
rect 462394 463818 462426 464054
rect 462662 463818 462746 464054
rect 462982 463818 463014 464054
rect 462394 463734 463014 463818
rect 462394 463498 462426 463734
rect 462662 463498 462746 463734
rect 462982 463498 463014 463734
rect 462394 430054 463014 463498
rect 462394 429818 462426 430054
rect 462662 429818 462746 430054
rect 462982 429818 463014 430054
rect 462394 429734 463014 429818
rect 462394 429498 462426 429734
rect 462662 429498 462746 429734
rect 462982 429498 463014 429734
rect 462394 396054 463014 429498
rect 462394 395818 462426 396054
rect 462662 395818 462746 396054
rect 462982 395818 463014 396054
rect 462394 395734 463014 395818
rect 462394 395498 462426 395734
rect 462662 395498 462746 395734
rect 462982 395498 463014 395734
rect 462394 362054 463014 395498
rect 462394 361818 462426 362054
rect 462662 361818 462746 362054
rect 462982 361818 463014 362054
rect 462394 361734 463014 361818
rect 462394 361498 462426 361734
rect 462662 361498 462746 361734
rect 462982 361498 463014 361734
rect 462394 328054 463014 361498
rect 462394 327818 462426 328054
rect 462662 327818 462746 328054
rect 462982 327818 463014 328054
rect 462394 327734 463014 327818
rect 462394 327498 462426 327734
rect 462662 327498 462746 327734
rect 462982 327498 463014 327734
rect 462394 294054 463014 327498
rect 462394 293818 462426 294054
rect 462662 293818 462746 294054
rect 462982 293818 463014 294054
rect 462394 293734 463014 293818
rect 462394 293498 462426 293734
rect 462662 293498 462746 293734
rect 462982 293498 463014 293734
rect 462394 260054 463014 293498
rect 462394 259818 462426 260054
rect 462662 259818 462746 260054
rect 462982 259818 463014 260054
rect 462394 259734 463014 259818
rect 462394 259498 462426 259734
rect 462662 259498 462746 259734
rect 462982 259498 463014 259734
rect 462394 226054 463014 259498
rect 462394 225818 462426 226054
rect 462662 225818 462746 226054
rect 462982 225818 463014 226054
rect 462394 225734 463014 225818
rect 462394 225498 462426 225734
rect 462662 225498 462746 225734
rect 462982 225498 463014 225734
rect 462394 192054 463014 225498
rect 462394 191818 462426 192054
rect 462662 191818 462746 192054
rect 462982 191818 463014 192054
rect 462394 191734 463014 191818
rect 462394 191498 462426 191734
rect 462662 191498 462746 191734
rect 462982 191498 463014 191734
rect 462394 158054 463014 191498
rect 462394 157818 462426 158054
rect 462662 157818 462746 158054
rect 462982 157818 463014 158054
rect 462394 157734 463014 157818
rect 462394 157498 462426 157734
rect 462662 157498 462746 157734
rect 462982 157498 463014 157734
rect 462394 124054 463014 157498
rect 462394 123818 462426 124054
rect 462662 123818 462746 124054
rect 462982 123818 463014 124054
rect 462394 123734 463014 123818
rect 462394 123498 462426 123734
rect 462662 123498 462746 123734
rect 462982 123498 463014 123734
rect 462394 90054 463014 123498
rect 462394 89818 462426 90054
rect 462662 89818 462746 90054
rect 462982 89818 463014 90054
rect 462394 89734 463014 89818
rect 462394 89498 462426 89734
rect 462662 89498 462746 89734
rect 462982 89498 463014 89734
rect 462394 56054 463014 89498
rect 462394 55818 462426 56054
rect 462662 55818 462746 56054
rect 462982 55818 463014 56054
rect 462394 55734 463014 55818
rect 462394 55498 462426 55734
rect 462662 55498 462746 55734
rect 462982 55498 463014 55734
rect 462394 22054 463014 55498
rect 462394 21818 462426 22054
rect 462662 21818 462746 22054
rect 462982 21818 463014 22054
rect 462394 21734 463014 21818
rect 462394 21498 462426 21734
rect 462662 21498 462746 21734
rect 462982 21498 463014 21734
rect 462394 -5146 463014 21498
rect 462394 -5382 462426 -5146
rect 462662 -5382 462746 -5146
rect 462982 -5382 463014 -5146
rect 462394 -5466 463014 -5382
rect 462394 -5702 462426 -5466
rect 462662 -5702 462746 -5466
rect 462982 -5702 463014 -5466
rect 462394 -7654 463014 -5702
rect 466114 710598 466734 711590
rect 466114 710362 466146 710598
rect 466382 710362 466466 710598
rect 466702 710362 466734 710598
rect 466114 710278 466734 710362
rect 466114 710042 466146 710278
rect 466382 710042 466466 710278
rect 466702 710042 466734 710278
rect 466114 671774 466734 710042
rect 466114 671538 466146 671774
rect 466382 671538 466466 671774
rect 466702 671538 466734 671774
rect 466114 671454 466734 671538
rect 466114 671218 466146 671454
rect 466382 671218 466466 671454
rect 466702 671218 466734 671454
rect 466114 637774 466734 671218
rect 466114 637538 466146 637774
rect 466382 637538 466466 637774
rect 466702 637538 466734 637774
rect 466114 637454 466734 637538
rect 466114 637218 466146 637454
rect 466382 637218 466466 637454
rect 466702 637218 466734 637454
rect 466114 603774 466734 637218
rect 466114 603538 466146 603774
rect 466382 603538 466466 603774
rect 466702 603538 466734 603774
rect 466114 603454 466734 603538
rect 466114 603218 466146 603454
rect 466382 603218 466466 603454
rect 466702 603218 466734 603454
rect 466114 569774 466734 603218
rect 466114 569538 466146 569774
rect 466382 569538 466466 569774
rect 466702 569538 466734 569774
rect 466114 569454 466734 569538
rect 466114 569218 466146 569454
rect 466382 569218 466466 569454
rect 466702 569218 466734 569454
rect 466114 535774 466734 569218
rect 466114 535538 466146 535774
rect 466382 535538 466466 535774
rect 466702 535538 466734 535774
rect 466114 535454 466734 535538
rect 466114 535218 466146 535454
rect 466382 535218 466466 535454
rect 466702 535218 466734 535454
rect 466114 501774 466734 535218
rect 466114 501538 466146 501774
rect 466382 501538 466466 501774
rect 466702 501538 466734 501774
rect 466114 501454 466734 501538
rect 466114 501218 466146 501454
rect 466382 501218 466466 501454
rect 466702 501218 466734 501454
rect 466114 467774 466734 501218
rect 466114 467538 466146 467774
rect 466382 467538 466466 467774
rect 466702 467538 466734 467774
rect 466114 467454 466734 467538
rect 466114 467218 466146 467454
rect 466382 467218 466466 467454
rect 466702 467218 466734 467454
rect 466114 433774 466734 467218
rect 466114 433538 466146 433774
rect 466382 433538 466466 433774
rect 466702 433538 466734 433774
rect 466114 433454 466734 433538
rect 466114 433218 466146 433454
rect 466382 433218 466466 433454
rect 466702 433218 466734 433454
rect 466114 399774 466734 433218
rect 466114 399538 466146 399774
rect 466382 399538 466466 399774
rect 466702 399538 466734 399774
rect 466114 399454 466734 399538
rect 466114 399218 466146 399454
rect 466382 399218 466466 399454
rect 466702 399218 466734 399454
rect 466114 365774 466734 399218
rect 466114 365538 466146 365774
rect 466382 365538 466466 365774
rect 466702 365538 466734 365774
rect 466114 365454 466734 365538
rect 466114 365218 466146 365454
rect 466382 365218 466466 365454
rect 466702 365218 466734 365454
rect 466114 331774 466734 365218
rect 466114 331538 466146 331774
rect 466382 331538 466466 331774
rect 466702 331538 466734 331774
rect 466114 331454 466734 331538
rect 466114 331218 466146 331454
rect 466382 331218 466466 331454
rect 466702 331218 466734 331454
rect 466114 297774 466734 331218
rect 466114 297538 466146 297774
rect 466382 297538 466466 297774
rect 466702 297538 466734 297774
rect 466114 297454 466734 297538
rect 466114 297218 466146 297454
rect 466382 297218 466466 297454
rect 466702 297218 466734 297454
rect 466114 263774 466734 297218
rect 466114 263538 466146 263774
rect 466382 263538 466466 263774
rect 466702 263538 466734 263774
rect 466114 263454 466734 263538
rect 466114 263218 466146 263454
rect 466382 263218 466466 263454
rect 466702 263218 466734 263454
rect 466114 229774 466734 263218
rect 466114 229538 466146 229774
rect 466382 229538 466466 229774
rect 466702 229538 466734 229774
rect 466114 229454 466734 229538
rect 466114 229218 466146 229454
rect 466382 229218 466466 229454
rect 466702 229218 466734 229454
rect 466114 195774 466734 229218
rect 466114 195538 466146 195774
rect 466382 195538 466466 195774
rect 466702 195538 466734 195774
rect 466114 195454 466734 195538
rect 466114 195218 466146 195454
rect 466382 195218 466466 195454
rect 466702 195218 466734 195454
rect 466114 161774 466734 195218
rect 466114 161538 466146 161774
rect 466382 161538 466466 161774
rect 466702 161538 466734 161774
rect 466114 161454 466734 161538
rect 466114 161218 466146 161454
rect 466382 161218 466466 161454
rect 466702 161218 466734 161454
rect 466114 127774 466734 161218
rect 466114 127538 466146 127774
rect 466382 127538 466466 127774
rect 466702 127538 466734 127774
rect 466114 127454 466734 127538
rect 466114 127218 466146 127454
rect 466382 127218 466466 127454
rect 466702 127218 466734 127454
rect 466114 93774 466734 127218
rect 466114 93538 466146 93774
rect 466382 93538 466466 93774
rect 466702 93538 466734 93774
rect 466114 93454 466734 93538
rect 466114 93218 466146 93454
rect 466382 93218 466466 93454
rect 466702 93218 466734 93454
rect 466114 59774 466734 93218
rect 466114 59538 466146 59774
rect 466382 59538 466466 59774
rect 466702 59538 466734 59774
rect 466114 59454 466734 59538
rect 466114 59218 466146 59454
rect 466382 59218 466466 59454
rect 466702 59218 466734 59454
rect 466114 25774 466734 59218
rect 466114 25538 466146 25774
rect 466382 25538 466466 25774
rect 466702 25538 466734 25774
rect 466114 25454 466734 25538
rect 466114 25218 466146 25454
rect 466382 25218 466466 25454
rect 466702 25218 466734 25454
rect 466114 -6106 466734 25218
rect 466114 -6342 466146 -6106
rect 466382 -6342 466466 -6106
rect 466702 -6342 466734 -6106
rect 466114 -6426 466734 -6342
rect 466114 -6662 466146 -6426
rect 466382 -6662 466466 -6426
rect 466702 -6662 466734 -6426
rect 466114 -7654 466734 -6662
rect 469834 711558 470454 711590
rect 469834 711322 469866 711558
rect 470102 711322 470186 711558
rect 470422 711322 470454 711558
rect 469834 711238 470454 711322
rect 469834 711002 469866 711238
rect 470102 711002 470186 711238
rect 470422 711002 470454 711238
rect 469834 675494 470454 711002
rect 469834 675258 469866 675494
rect 470102 675258 470186 675494
rect 470422 675258 470454 675494
rect 469834 675174 470454 675258
rect 469834 674938 469866 675174
rect 470102 674938 470186 675174
rect 470422 674938 470454 675174
rect 469834 641494 470454 674938
rect 469834 641258 469866 641494
rect 470102 641258 470186 641494
rect 470422 641258 470454 641494
rect 469834 641174 470454 641258
rect 469834 640938 469866 641174
rect 470102 640938 470186 641174
rect 470422 640938 470454 641174
rect 469834 607494 470454 640938
rect 469834 607258 469866 607494
rect 470102 607258 470186 607494
rect 470422 607258 470454 607494
rect 469834 607174 470454 607258
rect 469834 606938 469866 607174
rect 470102 606938 470186 607174
rect 470422 606938 470454 607174
rect 469834 573494 470454 606938
rect 469834 573258 469866 573494
rect 470102 573258 470186 573494
rect 470422 573258 470454 573494
rect 469834 573174 470454 573258
rect 469834 572938 469866 573174
rect 470102 572938 470186 573174
rect 470422 572938 470454 573174
rect 469834 539494 470454 572938
rect 469834 539258 469866 539494
rect 470102 539258 470186 539494
rect 470422 539258 470454 539494
rect 469834 539174 470454 539258
rect 469834 538938 469866 539174
rect 470102 538938 470186 539174
rect 470422 538938 470454 539174
rect 469834 505494 470454 538938
rect 469834 505258 469866 505494
rect 470102 505258 470186 505494
rect 470422 505258 470454 505494
rect 469834 505174 470454 505258
rect 469834 504938 469866 505174
rect 470102 504938 470186 505174
rect 470422 504938 470454 505174
rect 469834 471494 470454 504938
rect 469834 471258 469866 471494
rect 470102 471258 470186 471494
rect 470422 471258 470454 471494
rect 469834 471174 470454 471258
rect 469834 470938 469866 471174
rect 470102 470938 470186 471174
rect 470422 470938 470454 471174
rect 469834 437494 470454 470938
rect 469834 437258 469866 437494
rect 470102 437258 470186 437494
rect 470422 437258 470454 437494
rect 469834 437174 470454 437258
rect 469834 436938 469866 437174
rect 470102 436938 470186 437174
rect 470422 436938 470454 437174
rect 469834 403494 470454 436938
rect 469834 403258 469866 403494
rect 470102 403258 470186 403494
rect 470422 403258 470454 403494
rect 469834 403174 470454 403258
rect 469834 402938 469866 403174
rect 470102 402938 470186 403174
rect 470422 402938 470454 403174
rect 469834 369494 470454 402938
rect 469834 369258 469866 369494
rect 470102 369258 470186 369494
rect 470422 369258 470454 369494
rect 469834 369174 470454 369258
rect 469834 368938 469866 369174
rect 470102 368938 470186 369174
rect 470422 368938 470454 369174
rect 469834 335494 470454 368938
rect 469834 335258 469866 335494
rect 470102 335258 470186 335494
rect 470422 335258 470454 335494
rect 469834 335174 470454 335258
rect 469834 334938 469866 335174
rect 470102 334938 470186 335174
rect 470422 334938 470454 335174
rect 469834 301494 470454 334938
rect 469834 301258 469866 301494
rect 470102 301258 470186 301494
rect 470422 301258 470454 301494
rect 469834 301174 470454 301258
rect 469834 300938 469866 301174
rect 470102 300938 470186 301174
rect 470422 300938 470454 301174
rect 469834 267494 470454 300938
rect 469834 267258 469866 267494
rect 470102 267258 470186 267494
rect 470422 267258 470454 267494
rect 469834 267174 470454 267258
rect 469834 266938 469866 267174
rect 470102 266938 470186 267174
rect 470422 266938 470454 267174
rect 469834 233494 470454 266938
rect 469834 233258 469866 233494
rect 470102 233258 470186 233494
rect 470422 233258 470454 233494
rect 469834 233174 470454 233258
rect 469834 232938 469866 233174
rect 470102 232938 470186 233174
rect 470422 232938 470454 233174
rect 469834 199494 470454 232938
rect 469834 199258 469866 199494
rect 470102 199258 470186 199494
rect 470422 199258 470454 199494
rect 469834 199174 470454 199258
rect 469834 198938 469866 199174
rect 470102 198938 470186 199174
rect 470422 198938 470454 199174
rect 469834 165494 470454 198938
rect 469834 165258 469866 165494
rect 470102 165258 470186 165494
rect 470422 165258 470454 165494
rect 469834 165174 470454 165258
rect 469834 164938 469866 165174
rect 470102 164938 470186 165174
rect 470422 164938 470454 165174
rect 469834 131494 470454 164938
rect 469834 131258 469866 131494
rect 470102 131258 470186 131494
rect 470422 131258 470454 131494
rect 469834 131174 470454 131258
rect 469834 130938 469866 131174
rect 470102 130938 470186 131174
rect 470422 130938 470454 131174
rect 469834 97494 470454 130938
rect 469834 97258 469866 97494
rect 470102 97258 470186 97494
rect 470422 97258 470454 97494
rect 469834 97174 470454 97258
rect 469834 96938 469866 97174
rect 470102 96938 470186 97174
rect 470422 96938 470454 97174
rect 469834 63494 470454 96938
rect 469834 63258 469866 63494
rect 470102 63258 470186 63494
rect 470422 63258 470454 63494
rect 469834 63174 470454 63258
rect 469834 62938 469866 63174
rect 470102 62938 470186 63174
rect 470422 62938 470454 63174
rect 469834 29494 470454 62938
rect 469834 29258 469866 29494
rect 470102 29258 470186 29494
rect 470422 29258 470454 29494
rect 469834 29174 470454 29258
rect 469834 28938 469866 29174
rect 470102 28938 470186 29174
rect 470422 28938 470454 29174
rect 469834 -7066 470454 28938
rect 469834 -7302 469866 -7066
rect 470102 -7302 470186 -7066
rect 470422 -7302 470454 -7066
rect 469834 -7386 470454 -7302
rect 469834 -7622 469866 -7386
rect 470102 -7622 470186 -7386
rect 470422 -7622 470454 -7386
rect 469834 -7654 470454 -7622
rect 477794 704838 478414 711590
rect 477794 704602 477826 704838
rect 478062 704602 478146 704838
rect 478382 704602 478414 704838
rect 477794 704518 478414 704602
rect 477794 704282 477826 704518
rect 478062 704282 478146 704518
rect 478382 704282 478414 704518
rect 477794 683454 478414 704282
rect 477794 683218 477826 683454
rect 478062 683218 478146 683454
rect 478382 683218 478414 683454
rect 477794 683134 478414 683218
rect 477794 682898 477826 683134
rect 478062 682898 478146 683134
rect 478382 682898 478414 683134
rect 477794 649454 478414 682898
rect 477794 649218 477826 649454
rect 478062 649218 478146 649454
rect 478382 649218 478414 649454
rect 477794 649134 478414 649218
rect 477794 648898 477826 649134
rect 478062 648898 478146 649134
rect 478382 648898 478414 649134
rect 477794 615454 478414 648898
rect 477794 615218 477826 615454
rect 478062 615218 478146 615454
rect 478382 615218 478414 615454
rect 477794 615134 478414 615218
rect 477794 614898 477826 615134
rect 478062 614898 478146 615134
rect 478382 614898 478414 615134
rect 477794 581454 478414 614898
rect 477794 581218 477826 581454
rect 478062 581218 478146 581454
rect 478382 581218 478414 581454
rect 477794 581134 478414 581218
rect 477794 580898 477826 581134
rect 478062 580898 478146 581134
rect 478382 580898 478414 581134
rect 477794 547454 478414 580898
rect 477794 547218 477826 547454
rect 478062 547218 478146 547454
rect 478382 547218 478414 547454
rect 477794 547134 478414 547218
rect 477794 546898 477826 547134
rect 478062 546898 478146 547134
rect 478382 546898 478414 547134
rect 477794 513454 478414 546898
rect 477794 513218 477826 513454
rect 478062 513218 478146 513454
rect 478382 513218 478414 513454
rect 477794 513134 478414 513218
rect 477794 512898 477826 513134
rect 478062 512898 478146 513134
rect 478382 512898 478414 513134
rect 477794 479454 478414 512898
rect 477794 479218 477826 479454
rect 478062 479218 478146 479454
rect 478382 479218 478414 479454
rect 477794 479134 478414 479218
rect 477794 478898 477826 479134
rect 478062 478898 478146 479134
rect 478382 478898 478414 479134
rect 477794 445454 478414 478898
rect 477794 445218 477826 445454
rect 478062 445218 478146 445454
rect 478382 445218 478414 445454
rect 477794 445134 478414 445218
rect 477794 444898 477826 445134
rect 478062 444898 478146 445134
rect 478382 444898 478414 445134
rect 477794 411454 478414 444898
rect 477794 411218 477826 411454
rect 478062 411218 478146 411454
rect 478382 411218 478414 411454
rect 477794 411134 478414 411218
rect 477794 410898 477826 411134
rect 478062 410898 478146 411134
rect 478382 410898 478414 411134
rect 477794 377454 478414 410898
rect 477794 377218 477826 377454
rect 478062 377218 478146 377454
rect 478382 377218 478414 377454
rect 477794 377134 478414 377218
rect 477794 376898 477826 377134
rect 478062 376898 478146 377134
rect 478382 376898 478414 377134
rect 477794 343454 478414 376898
rect 477794 343218 477826 343454
rect 478062 343218 478146 343454
rect 478382 343218 478414 343454
rect 477794 343134 478414 343218
rect 477794 342898 477826 343134
rect 478062 342898 478146 343134
rect 478382 342898 478414 343134
rect 477794 309454 478414 342898
rect 477794 309218 477826 309454
rect 478062 309218 478146 309454
rect 478382 309218 478414 309454
rect 477794 309134 478414 309218
rect 477794 308898 477826 309134
rect 478062 308898 478146 309134
rect 478382 308898 478414 309134
rect 477794 275454 478414 308898
rect 477794 275218 477826 275454
rect 478062 275218 478146 275454
rect 478382 275218 478414 275454
rect 477794 275134 478414 275218
rect 477794 274898 477826 275134
rect 478062 274898 478146 275134
rect 478382 274898 478414 275134
rect 477794 241454 478414 274898
rect 477794 241218 477826 241454
rect 478062 241218 478146 241454
rect 478382 241218 478414 241454
rect 477794 241134 478414 241218
rect 477794 240898 477826 241134
rect 478062 240898 478146 241134
rect 478382 240898 478414 241134
rect 477794 207454 478414 240898
rect 477794 207218 477826 207454
rect 478062 207218 478146 207454
rect 478382 207218 478414 207454
rect 477794 207134 478414 207218
rect 477794 206898 477826 207134
rect 478062 206898 478146 207134
rect 478382 206898 478414 207134
rect 477794 173454 478414 206898
rect 477794 173218 477826 173454
rect 478062 173218 478146 173454
rect 478382 173218 478414 173454
rect 477794 173134 478414 173218
rect 477794 172898 477826 173134
rect 478062 172898 478146 173134
rect 478382 172898 478414 173134
rect 477794 139454 478414 172898
rect 477794 139218 477826 139454
rect 478062 139218 478146 139454
rect 478382 139218 478414 139454
rect 477794 139134 478414 139218
rect 477794 138898 477826 139134
rect 478062 138898 478146 139134
rect 478382 138898 478414 139134
rect 477794 105454 478414 138898
rect 477794 105218 477826 105454
rect 478062 105218 478146 105454
rect 478382 105218 478414 105454
rect 477794 105134 478414 105218
rect 477794 104898 477826 105134
rect 478062 104898 478146 105134
rect 478382 104898 478414 105134
rect 477794 71454 478414 104898
rect 477794 71218 477826 71454
rect 478062 71218 478146 71454
rect 478382 71218 478414 71454
rect 477794 71134 478414 71218
rect 477794 70898 477826 71134
rect 478062 70898 478146 71134
rect 478382 70898 478414 71134
rect 477794 37454 478414 70898
rect 477794 37218 477826 37454
rect 478062 37218 478146 37454
rect 478382 37218 478414 37454
rect 477794 37134 478414 37218
rect 477794 36898 477826 37134
rect 478062 36898 478146 37134
rect 478382 36898 478414 37134
rect 477794 3454 478414 36898
rect 477794 3218 477826 3454
rect 478062 3218 478146 3454
rect 478382 3218 478414 3454
rect 477794 3134 478414 3218
rect 477794 2898 477826 3134
rect 478062 2898 478146 3134
rect 478382 2898 478414 3134
rect 477794 -346 478414 2898
rect 477794 -582 477826 -346
rect 478062 -582 478146 -346
rect 478382 -582 478414 -346
rect 477794 -666 478414 -582
rect 477794 -902 477826 -666
rect 478062 -902 478146 -666
rect 478382 -902 478414 -666
rect 477794 -7654 478414 -902
rect 481514 705798 482134 711590
rect 481514 705562 481546 705798
rect 481782 705562 481866 705798
rect 482102 705562 482134 705798
rect 481514 705478 482134 705562
rect 481514 705242 481546 705478
rect 481782 705242 481866 705478
rect 482102 705242 482134 705478
rect 481514 687174 482134 705242
rect 481514 686938 481546 687174
rect 481782 686938 481866 687174
rect 482102 686938 482134 687174
rect 481514 686854 482134 686938
rect 481514 686618 481546 686854
rect 481782 686618 481866 686854
rect 482102 686618 482134 686854
rect 481514 653174 482134 686618
rect 481514 652938 481546 653174
rect 481782 652938 481866 653174
rect 482102 652938 482134 653174
rect 481514 652854 482134 652938
rect 481514 652618 481546 652854
rect 481782 652618 481866 652854
rect 482102 652618 482134 652854
rect 481514 619174 482134 652618
rect 481514 618938 481546 619174
rect 481782 618938 481866 619174
rect 482102 618938 482134 619174
rect 481514 618854 482134 618938
rect 481514 618618 481546 618854
rect 481782 618618 481866 618854
rect 482102 618618 482134 618854
rect 481514 585174 482134 618618
rect 481514 584938 481546 585174
rect 481782 584938 481866 585174
rect 482102 584938 482134 585174
rect 481514 584854 482134 584938
rect 481514 584618 481546 584854
rect 481782 584618 481866 584854
rect 482102 584618 482134 584854
rect 481514 551174 482134 584618
rect 481514 550938 481546 551174
rect 481782 550938 481866 551174
rect 482102 550938 482134 551174
rect 481514 550854 482134 550938
rect 481514 550618 481546 550854
rect 481782 550618 481866 550854
rect 482102 550618 482134 550854
rect 481514 517174 482134 550618
rect 481514 516938 481546 517174
rect 481782 516938 481866 517174
rect 482102 516938 482134 517174
rect 481514 516854 482134 516938
rect 481514 516618 481546 516854
rect 481782 516618 481866 516854
rect 482102 516618 482134 516854
rect 481514 483174 482134 516618
rect 481514 482938 481546 483174
rect 481782 482938 481866 483174
rect 482102 482938 482134 483174
rect 481514 482854 482134 482938
rect 481514 482618 481546 482854
rect 481782 482618 481866 482854
rect 482102 482618 482134 482854
rect 481514 449174 482134 482618
rect 481514 448938 481546 449174
rect 481782 448938 481866 449174
rect 482102 448938 482134 449174
rect 481514 448854 482134 448938
rect 481514 448618 481546 448854
rect 481782 448618 481866 448854
rect 482102 448618 482134 448854
rect 481514 415174 482134 448618
rect 481514 414938 481546 415174
rect 481782 414938 481866 415174
rect 482102 414938 482134 415174
rect 481514 414854 482134 414938
rect 481514 414618 481546 414854
rect 481782 414618 481866 414854
rect 482102 414618 482134 414854
rect 481514 381174 482134 414618
rect 481514 380938 481546 381174
rect 481782 380938 481866 381174
rect 482102 380938 482134 381174
rect 481514 380854 482134 380938
rect 481514 380618 481546 380854
rect 481782 380618 481866 380854
rect 482102 380618 482134 380854
rect 481514 347174 482134 380618
rect 481514 346938 481546 347174
rect 481782 346938 481866 347174
rect 482102 346938 482134 347174
rect 481514 346854 482134 346938
rect 481514 346618 481546 346854
rect 481782 346618 481866 346854
rect 482102 346618 482134 346854
rect 481514 313174 482134 346618
rect 481514 312938 481546 313174
rect 481782 312938 481866 313174
rect 482102 312938 482134 313174
rect 481514 312854 482134 312938
rect 481514 312618 481546 312854
rect 481782 312618 481866 312854
rect 482102 312618 482134 312854
rect 481514 279174 482134 312618
rect 481514 278938 481546 279174
rect 481782 278938 481866 279174
rect 482102 278938 482134 279174
rect 481514 278854 482134 278938
rect 481514 278618 481546 278854
rect 481782 278618 481866 278854
rect 482102 278618 482134 278854
rect 481514 245174 482134 278618
rect 481514 244938 481546 245174
rect 481782 244938 481866 245174
rect 482102 244938 482134 245174
rect 481514 244854 482134 244938
rect 481514 244618 481546 244854
rect 481782 244618 481866 244854
rect 482102 244618 482134 244854
rect 481514 211174 482134 244618
rect 481514 210938 481546 211174
rect 481782 210938 481866 211174
rect 482102 210938 482134 211174
rect 481514 210854 482134 210938
rect 481514 210618 481546 210854
rect 481782 210618 481866 210854
rect 482102 210618 482134 210854
rect 481514 177174 482134 210618
rect 481514 176938 481546 177174
rect 481782 176938 481866 177174
rect 482102 176938 482134 177174
rect 481514 176854 482134 176938
rect 481514 176618 481546 176854
rect 481782 176618 481866 176854
rect 482102 176618 482134 176854
rect 481514 143174 482134 176618
rect 481514 142938 481546 143174
rect 481782 142938 481866 143174
rect 482102 142938 482134 143174
rect 481514 142854 482134 142938
rect 481514 142618 481546 142854
rect 481782 142618 481866 142854
rect 482102 142618 482134 142854
rect 481514 109174 482134 142618
rect 481514 108938 481546 109174
rect 481782 108938 481866 109174
rect 482102 108938 482134 109174
rect 481514 108854 482134 108938
rect 481514 108618 481546 108854
rect 481782 108618 481866 108854
rect 482102 108618 482134 108854
rect 481514 75174 482134 108618
rect 481514 74938 481546 75174
rect 481782 74938 481866 75174
rect 482102 74938 482134 75174
rect 481514 74854 482134 74938
rect 481514 74618 481546 74854
rect 481782 74618 481866 74854
rect 482102 74618 482134 74854
rect 481514 41174 482134 74618
rect 481514 40938 481546 41174
rect 481782 40938 481866 41174
rect 482102 40938 482134 41174
rect 481514 40854 482134 40938
rect 481514 40618 481546 40854
rect 481782 40618 481866 40854
rect 482102 40618 482134 40854
rect 481514 7174 482134 40618
rect 481514 6938 481546 7174
rect 481782 6938 481866 7174
rect 482102 6938 482134 7174
rect 481514 6854 482134 6938
rect 481514 6618 481546 6854
rect 481782 6618 481866 6854
rect 482102 6618 482134 6854
rect 481514 -1306 482134 6618
rect 481514 -1542 481546 -1306
rect 481782 -1542 481866 -1306
rect 482102 -1542 482134 -1306
rect 481514 -1626 482134 -1542
rect 481514 -1862 481546 -1626
rect 481782 -1862 481866 -1626
rect 482102 -1862 482134 -1626
rect 481514 -7654 482134 -1862
rect 485234 706758 485854 711590
rect 485234 706522 485266 706758
rect 485502 706522 485586 706758
rect 485822 706522 485854 706758
rect 485234 706438 485854 706522
rect 485234 706202 485266 706438
rect 485502 706202 485586 706438
rect 485822 706202 485854 706438
rect 485234 690894 485854 706202
rect 485234 690658 485266 690894
rect 485502 690658 485586 690894
rect 485822 690658 485854 690894
rect 485234 690574 485854 690658
rect 485234 690338 485266 690574
rect 485502 690338 485586 690574
rect 485822 690338 485854 690574
rect 485234 656894 485854 690338
rect 485234 656658 485266 656894
rect 485502 656658 485586 656894
rect 485822 656658 485854 656894
rect 485234 656574 485854 656658
rect 485234 656338 485266 656574
rect 485502 656338 485586 656574
rect 485822 656338 485854 656574
rect 485234 622894 485854 656338
rect 485234 622658 485266 622894
rect 485502 622658 485586 622894
rect 485822 622658 485854 622894
rect 485234 622574 485854 622658
rect 485234 622338 485266 622574
rect 485502 622338 485586 622574
rect 485822 622338 485854 622574
rect 485234 588894 485854 622338
rect 485234 588658 485266 588894
rect 485502 588658 485586 588894
rect 485822 588658 485854 588894
rect 485234 588574 485854 588658
rect 485234 588338 485266 588574
rect 485502 588338 485586 588574
rect 485822 588338 485854 588574
rect 485234 554894 485854 588338
rect 485234 554658 485266 554894
rect 485502 554658 485586 554894
rect 485822 554658 485854 554894
rect 485234 554574 485854 554658
rect 485234 554338 485266 554574
rect 485502 554338 485586 554574
rect 485822 554338 485854 554574
rect 485234 520894 485854 554338
rect 485234 520658 485266 520894
rect 485502 520658 485586 520894
rect 485822 520658 485854 520894
rect 485234 520574 485854 520658
rect 485234 520338 485266 520574
rect 485502 520338 485586 520574
rect 485822 520338 485854 520574
rect 485234 486894 485854 520338
rect 485234 486658 485266 486894
rect 485502 486658 485586 486894
rect 485822 486658 485854 486894
rect 485234 486574 485854 486658
rect 485234 486338 485266 486574
rect 485502 486338 485586 486574
rect 485822 486338 485854 486574
rect 485234 452894 485854 486338
rect 485234 452658 485266 452894
rect 485502 452658 485586 452894
rect 485822 452658 485854 452894
rect 485234 452574 485854 452658
rect 485234 452338 485266 452574
rect 485502 452338 485586 452574
rect 485822 452338 485854 452574
rect 485234 418894 485854 452338
rect 485234 418658 485266 418894
rect 485502 418658 485586 418894
rect 485822 418658 485854 418894
rect 485234 418574 485854 418658
rect 485234 418338 485266 418574
rect 485502 418338 485586 418574
rect 485822 418338 485854 418574
rect 485234 384894 485854 418338
rect 485234 384658 485266 384894
rect 485502 384658 485586 384894
rect 485822 384658 485854 384894
rect 485234 384574 485854 384658
rect 485234 384338 485266 384574
rect 485502 384338 485586 384574
rect 485822 384338 485854 384574
rect 485234 350894 485854 384338
rect 485234 350658 485266 350894
rect 485502 350658 485586 350894
rect 485822 350658 485854 350894
rect 485234 350574 485854 350658
rect 485234 350338 485266 350574
rect 485502 350338 485586 350574
rect 485822 350338 485854 350574
rect 485234 316894 485854 350338
rect 485234 316658 485266 316894
rect 485502 316658 485586 316894
rect 485822 316658 485854 316894
rect 485234 316574 485854 316658
rect 485234 316338 485266 316574
rect 485502 316338 485586 316574
rect 485822 316338 485854 316574
rect 485234 282894 485854 316338
rect 485234 282658 485266 282894
rect 485502 282658 485586 282894
rect 485822 282658 485854 282894
rect 485234 282574 485854 282658
rect 485234 282338 485266 282574
rect 485502 282338 485586 282574
rect 485822 282338 485854 282574
rect 485234 248894 485854 282338
rect 485234 248658 485266 248894
rect 485502 248658 485586 248894
rect 485822 248658 485854 248894
rect 485234 248574 485854 248658
rect 485234 248338 485266 248574
rect 485502 248338 485586 248574
rect 485822 248338 485854 248574
rect 485234 214894 485854 248338
rect 485234 214658 485266 214894
rect 485502 214658 485586 214894
rect 485822 214658 485854 214894
rect 485234 214574 485854 214658
rect 485234 214338 485266 214574
rect 485502 214338 485586 214574
rect 485822 214338 485854 214574
rect 485234 180894 485854 214338
rect 485234 180658 485266 180894
rect 485502 180658 485586 180894
rect 485822 180658 485854 180894
rect 485234 180574 485854 180658
rect 485234 180338 485266 180574
rect 485502 180338 485586 180574
rect 485822 180338 485854 180574
rect 485234 146894 485854 180338
rect 485234 146658 485266 146894
rect 485502 146658 485586 146894
rect 485822 146658 485854 146894
rect 485234 146574 485854 146658
rect 485234 146338 485266 146574
rect 485502 146338 485586 146574
rect 485822 146338 485854 146574
rect 485234 112894 485854 146338
rect 485234 112658 485266 112894
rect 485502 112658 485586 112894
rect 485822 112658 485854 112894
rect 485234 112574 485854 112658
rect 485234 112338 485266 112574
rect 485502 112338 485586 112574
rect 485822 112338 485854 112574
rect 485234 78894 485854 112338
rect 485234 78658 485266 78894
rect 485502 78658 485586 78894
rect 485822 78658 485854 78894
rect 485234 78574 485854 78658
rect 485234 78338 485266 78574
rect 485502 78338 485586 78574
rect 485822 78338 485854 78574
rect 485234 44894 485854 78338
rect 485234 44658 485266 44894
rect 485502 44658 485586 44894
rect 485822 44658 485854 44894
rect 485234 44574 485854 44658
rect 485234 44338 485266 44574
rect 485502 44338 485586 44574
rect 485822 44338 485854 44574
rect 485234 10894 485854 44338
rect 485234 10658 485266 10894
rect 485502 10658 485586 10894
rect 485822 10658 485854 10894
rect 485234 10574 485854 10658
rect 485234 10338 485266 10574
rect 485502 10338 485586 10574
rect 485822 10338 485854 10574
rect 485234 -2266 485854 10338
rect 485234 -2502 485266 -2266
rect 485502 -2502 485586 -2266
rect 485822 -2502 485854 -2266
rect 485234 -2586 485854 -2502
rect 485234 -2822 485266 -2586
rect 485502 -2822 485586 -2586
rect 485822 -2822 485854 -2586
rect 485234 -7654 485854 -2822
rect 488954 707718 489574 711590
rect 488954 707482 488986 707718
rect 489222 707482 489306 707718
rect 489542 707482 489574 707718
rect 488954 707398 489574 707482
rect 488954 707162 488986 707398
rect 489222 707162 489306 707398
rect 489542 707162 489574 707398
rect 488954 694614 489574 707162
rect 488954 694378 488986 694614
rect 489222 694378 489306 694614
rect 489542 694378 489574 694614
rect 488954 694294 489574 694378
rect 488954 694058 488986 694294
rect 489222 694058 489306 694294
rect 489542 694058 489574 694294
rect 488954 660614 489574 694058
rect 488954 660378 488986 660614
rect 489222 660378 489306 660614
rect 489542 660378 489574 660614
rect 488954 660294 489574 660378
rect 488954 660058 488986 660294
rect 489222 660058 489306 660294
rect 489542 660058 489574 660294
rect 488954 626614 489574 660058
rect 488954 626378 488986 626614
rect 489222 626378 489306 626614
rect 489542 626378 489574 626614
rect 488954 626294 489574 626378
rect 488954 626058 488986 626294
rect 489222 626058 489306 626294
rect 489542 626058 489574 626294
rect 488954 592614 489574 626058
rect 488954 592378 488986 592614
rect 489222 592378 489306 592614
rect 489542 592378 489574 592614
rect 488954 592294 489574 592378
rect 488954 592058 488986 592294
rect 489222 592058 489306 592294
rect 489542 592058 489574 592294
rect 488954 558614 489574 592058
rect 488954 558378 488986 558614
rect 489222 558378 489306 558614
rect 489542 558378 489574 558614
rect 488954 558294 489574 558378
rect 488954 558058 488986 558294
rect 489222 558058 489306 558294
rect 489542 558058 489574 558294
rect 488954 524614 489574 558058
rect 488954 524378 488986 524614
rect 489222 524378 489306 524614
rect 489542 524378 489574 524614
rect 488954 524294 489574 524378
rect 488954 524058 488986 524294
rect 489222 524058 489306 524294
rect 489542 524058 489574 524294
rect 488954 490614 489574 524058
rect 488954 490378 488986 490614
rect 489222 490378 489306 490614
rect 489542 490378 489574 490614
rect 488954 490294 489574 490378
rect 488954 490058 488986 490294
rect 489222 490058 489306 490294
rect 489542 490058 489574 490294
rect 488954 456614 489574 490058
rect 488954 456378 488986 456614
rect 489222 456378 489306 456614
rect 489542 456378 489574 456614
rect 488954 456294 489574 456378
rect 488954 456058 488986 456294
rect 489222 456058 489306 456294
rect 489542 456058 489574 456294
rect 488954 422614 489574 456058
rect 488954 422378 488986 422614
rect 489222 422378 489306 422614
rect 489542 422378 489574 422614
rect 488954 422294 489574 422378
rect 488954 422058 488986 422294
rect 489222 422058 489306 422294
rect 489542 422058 489574 422294
rect 488954 388614 489574 422058
rect 488954 388378 488986 388614
rect 489222 388378 489306 388614
rect 489542 388378 489574 388614
rect 488954 388294 489574 388378
rect 488954 388058 488986 388294
rect 489222 388058 489306 388294
rect 489542 388058 489574 388294
rect 488954 354614 489574 388058
rect 488954 354378 488986 354614
rect 489222 354378 489306 354614
rect 489542 354378 489574 354614
rect 488954 354294 489574 354378
rect 488954 354058 488986 354294
rect 489222 354058 489306 354294
rect 489542 354058 489574 354294
rect 488954 320614 489574 354058
rect 488954 320378 488986 320614
rect 489222 320378 489306 320614
rect 489542 320378 489574 320614
rect 488954 320294 489574 320378
rect 488954 320058 488986 320294
rect 489222 320058 489306 320294
rect 489542 320058 489574 320294
rect 488954 286614 489574 320058
rect 488954 286378 488986 286614
rect 489222 286378 489306 286614
rect 489542 286378 489574 286614
rect 488954 286294 489574 286378
rect 488954 286058 488986 286294
rect 489222 286058 489306 286294
rect 489542 286058 489574 286294
rect 488954 252614 489574 286058
rect 488954 252378 488986 252614
rect 489222 252378 489306 252614
rect 489542 252378 489574 252614
rect 488954 252294 489574 252378
rect 488954 252058 488986 252294
rect 489222 252058 489306 252294
rect 489542 252058 489574 252294
rect 488954 218614 489574 252058
rect 488954 218378 488986 218614
rect 489222 218378 489306 218614
rect 489542 218378 489574 218614
rect 488954 218294 489574 218378
rect 488954 218058 488986 218294
rect 489222 218058 489306 218294
rect 489542 218058 489574 218294
rect 488954 184614 489574 218058
rect 488954 184378 488986 184614
rect 489222 184378 489306 184614
rect 489542 184378 489574 184614
rect 488954 184294 489574 184378
rect 488954 184058 488986 184294
rect 489222 184058 489306 184294
rect 489542 184058 489574 184294
rect 488954 150614 489574 184058
rect 488954 150378 488986 150614
rect 489222 150378 489306 150614
rect 489542 150378 489574 150614
rect 488954 150294 489574 150378
rect 488954 150058 488986 150294
rect 489222 150058 489306 150294
rect 489542 150058 489574 150294
rect 488954 116614 489574 150058
rect 488954 116378 488986 116614
rect 489222 116378 489306 116614
rect 489542 116378 489574 116614
rect 488954 116294 489574 116378
rect 488954 116058 488986 116294
rect 489222 116058 489306 116294
rect 489542 116058 489574 116294
rect 488954 82614 489574 116058
rect 488954 82378 488986 82614
rect 489222 82378 489306 82614
rect 489542 82378 489574 82614
rect 488954 82294 489574 82378
rect 488954 82058 488986 82294
rect 489222 82058 489306 82294
rect 489542 82058 489574 82294
rect 488954 48614 489574 82058
rect 488954 48378 488986 48614
rect 489222 48378 489306 48614
rect 489542 48378 489574 48614
rect 488954 48294 489574 48378
rect 488954 48058 488986 48294
rect 489222 48058 489306 48294
rect 489542 48058 489574 48294
rect 488954 14614 489574 48058
rect 488954 14378 488986 14614
rect 489222 14378 489306 14614
rect 489542 14378 489574 14614
rect 488954 14294 489574 14378
rect 488954 14058 488986 14294
rect 489222 14058 489306 14294
rect 489542 14058 489574 14294
rect 488954 -3226 489574 14058
rect 488954 -3462 488986 -3226
rect 489222 -3462 489306 -3226
rect 489542 -3462 489574 -3226
rect 488954 -3546 489574 -3462
rect 488954 -3782 488986 -3546
rect 489222 -3782 489306 -3546
rect 489542 -3782 489574 -3546
rect 488954 -7654 489574 -3782
rect 492674 708678 493294 711590
rect 492674 708442 492706 708678
rect 492942 708442 493026 708678
rect 493262 708442 493294 708678
rect 492674 708358 493294 708442
rect 492674 708122 492706 708358
rect 492942 708122 493026 708358
rect 493262 708122 493294 708358
rect 492674 698334 493294 708122
rect 492674 698098 492706 698334
rect 492942 698098 493026 698334
rect 493262 698098 493294 698334
rect 492674 698014 493294 698098
rect 492674 697778 492706 698014
rect 492942 697778 493026 698014
rect 493262 697778 493294 698014
rect 492674 664334 493294 697778
rect 492674 664098 492706 664334
rect 492942 664098 493026 664334
rect 493262 664098 493294 664334
rect 492674 664014 493294 664098
rect 492674 663778 492706 664014
rect 492942 663778 493026 664014
rect 493262 663778 493294 664014
rect 492674 630334 493294 663778
rect 492674 630098 492706 630334
rect 492942 630098 493026 630334
rect 493262 630098 493294 630334
rect 492674 630014 493294 630098
rect 492674 629778 492706 630014
rect 492942 629778 493026 630014
rect 493262 629778 493294 630014
rect 492674 596334 493294 629778
rect 492674 596098 492706 596334
rect 492942 596098 493026 596334
rect 493262 596098 493294 596334
rect 492674 596014 493294 596098
rect 492674 595778 492706 596014
rect 492942 595778 493026 596014
rect 493262 595778 493294 596014
rect 492674 562334 493294 595778
rect 492674 562098 492706 562334
rect 492942 562098 493026 562334
rect 493262 562098 493294 562334
rect 492674 562014 493294 562098
rect 492674 561778 492706 562014
rect 492942 561778 493026 562014
rect 493262 561778 493294 562014
rect 492674 528334 493294 561778
rect 492674 528098 492706 528334
rect 492942 528098 493026 528334
rect 493262 528098 493294 528334
rect 492674 528014 493294 528098
rect 492674 527778 492706 528014
rect 492942 527778 493026 528014
rect 493262 527778 493294 528014
rect 492674 494334 493294 527778
rect 492674 494098 492706 494334
rect 492942 494098 493026 494334
rect 493262 494098 493294 494334
rect 492674 494014 493294 494098
rect 492674 493778 492706 494014
rect 492942 493778 493026 494014
rect 493262 493778 493294 494014
rect 492674 460334 493294 493778
rect 492674 460098 492706 460334
rect 492942 460098 493026 460334
rect 493262 460098 493294 460334
rect 492674 460014 493294 460098
rect 492674 459778 492706 460014
rect 492942 459778 493026 460014
rect 493262 459778 493294 460014
rect 492674 426334 493294 459778
rect 492674 426098 492706 426334
rect 492942 426098 493026 426334
rect 493262 426098 493294 426334
rect 492674 426014 493294 426098
rect 492674 425778 492706 426014
rect 492942 425778 493026 426014
rect 493262 425778 493294 426014
rect 492674 392334 493294 425778
rect 492674 392098 492706 392334
rect 492942 392098 493026 392334
rect 493262 392098 493294 392334
rect 492674 392014 493294 392098
rect 492674 391778 492706 392014
rect 492942 391778 493026 392014
rect 493262 391778 493294 392014
rect 492674 358334 493294 391778
rect 492674 358098 492706 358334
rect 492942 358098 493026 358334
rect 493262 358098 493294 358334
rect 492674 358014 493294 358098
rect 492674 357778 492706 358014
rect 492942 357778 493026 358014
rect 493262 357778 493294 358014
rect 492674 324334 493294 357778
rect 492674 324098 492706 324334
rect 492942 324098 493026 324334
rect 493262 324098 493294 324334
rect 492674 324014 493294 324098
rect 492674 323778 492706 324014
rect 492942 323778 493026 324014
rect 493262 323778 493294 324014
rect 492674 290334 493294 323778
rect 492674 290098 492706 290334
rect 492942 290098 493026 290334
rect 493262 290098 493294 290334
rect 492674 290014 493294 290098
rect 492674 289778 492706 290014
rect 492942 289778 493026 290014
rect 493262 289778 493294 290014
rect 492674 256334 493294 289778
rect 492674 256098 492706 256334
rect 492942 256098 493026 256334
rect 493262 256098 493294 256334
rect 492674 256014 493294 256098
rect 492674 255778 492706 256014
rect 492942 255778 493026 256014
rect 493262 255778 493294 256014
rect 492674 222334 493294 255778
rect 492674 222098 492706 222334
rect 492942 222098 493026 222334
rect 493262 222098 493294 222334
rect 492674 222014 493294 222098
rect 492674 221778 492706 222014
rect 492942 221778 493026 222014
rect 493262 221778 493294 222014
rect 492674 188334 493294 221778
rect 492674 188098 492706 188334
rect 492942 188098 493026 188334
rect 493262 188098 493294 188334
rect 492674 188014 493294 188098
rect 492674 187778 492706 188014
rect 492942 187778 493026 188014
rect 493262 187778 493294 188014
rect 492674 154334 493294 187778
rect 492674 154098 492706 154334
rect 492942 154098 493026 154334
rect 493262 154098 493294 154334
rect 492674 154014 493294 154098
rect 492674 153778 492706 154014
rect 492942 153778 493026 154014
rect 493262 153778 493294 154014
rect 492674 120334 493294 153778
rect 492674 120098 492706 120334
rect 492942 120098 493026 120334
rect 493262 120098 493294 120334
rect 492674 120014 493294 120098
rect 492674 119778 492706 120014
rect 492942 119778 493026 120014
rect 493262 119778 493294 120014
rect 492674 86334 493294 119778
rect 492674 86098 492706 86334
rect 492942 86098 493026 86334
rect 493262 86098 493294 86334
rect 492674 86014 493294 86098
rect 492674 85778 492706 86014
rect 492942 85778 493026 86014
rect 493262 85778 493294 86014
rect 492674 52334 493294 85778
rect 492674 52098 492706 52334
rect 492942 52098 493026 52334
rect 493262 52098 493294 52334
rect 492674 52014 493294 52098
rect 492674 51778 492706 52014
rect 492942 51778 493026 52014
rect 493262 51778 493294 52014
rect 492674 18334 493294 51778
rect 492674 18098 492706 18334
rect 492942 18098 493026 18334
rect 493262 18098 493294 18334
rect 492674 18014 493294 18098
rect 492674 17778 492706 18014
rect 492942 17778 493026 18014
rect 493262 17778 493294 18014
rect 492674 -4186 493294 17778
rect 492674 -4422 492706 -4186
rect 492942 -4422 493026 -4186
rect 493262 -4422 493294 -4186
rect 492674 -4506 493294 -4422
rect 492674 -4742 492706 -4506
rect 492942 -4742 493026 -4506
rect 493262 -4742 493294 -4506
rect 492674 -7654 493294 -4742
rect 496394 709638 497014 711590
rect 496394 709402 496426 709638
rect 496662 709402 496746 709638
rect 496982 709402 497014 709638
rect 496394 709318 497014 709402
rect 496394 709082 496426 709318
rect 496662 709082 496746 709318
rect 496982 709082 497014 709318
rect 496394 668054 497014 709082
rect 496394 667818 496426 668054
rect 496662 667818 496746 668054
rect 496982 667818 497014 668054
rect 496394 667734 497014 667818
rect 496394 667498 496426 667734
rect 496662 667498 496746 667734
rect 496982 667498 497014 667734
rect 496394 634054 497014 667498
rect 496394 633818 496426 634054
rect 496662 633818 496746 634054
rect 496982 633818 497014 634054
rect 496394 633734 497014 633818
rect 496394 633498 496426 633734
rect 496662 633498 496746 633734
rect 496982 633498 497014 633734
rect 496394 600054 497014 633498
rect 496394 599818 496426 600054
rect 496662 599818 496746 600054
rect 496982 599818 497014 600054
rect 496394 599734 497014 599818
rect 496394 599498 496426 599734
rect 496662 599498 496746 599734
rect 496982 599498 497014 599734
rect 496394 566054 497014 599498
rect 496394 565818 496426 566054
rect 496662 565818 496746 566054
rect 496982 565818 497014 566054
rect 496394 565734 497014 565818
rect 496394 565498 496426 565734
rect 496662 565498 496746 565734
rect 496982 565498 497014 565734
rect 496394 532054 497014 565498
rect 496394 531818 496426 532054
rect 496662 531818 496746 532054
rect 496982 531818 497014 532054
rect 496394 531734 497014 531818
rect 496394 531498 496426 531734
rect 496662 531498 496746 531734
rect 496982 531498 497014 531734
rect 496394 498054 497014 531498
rect 496394 497818 496426 498054
rect 496662 497818 496746 498054
rect 496982 497818 497014 498054
rect 496394 497734 497014 497818
rect 496394 497498 496426 497734
rect 496662 497498 496746 497734
rect 496982 497498 497014 497734
rect 496394 464054 497014 497498
rect 496394 463818 496426 464054
rect 496662 463818 496746 464054
rect 496982 463818 497014 464054
rect 496394 463734 497014 463818
rect 496394 463498 496426 463734
rect 496662 463498 496746 463734
rect 496982 463498 497014 463734
rect 496394 430054 497014 463498
rect 496394 429818 496426 430054
rect 496662 429818 496746 430054
rect 496982 429818 497014 430054
rect 496394 429734 497014 429818
rect 496394 429498 496426 429734
rect 496662 429498 496746 429734
rect 496982 429498 497014 429734
rect 496394 396054 497014 429498
rect 496394 395818 496426 396054
rect 496662 395818 496746 396054
rect 496982 395818 497014 396054
rect 496394 395734 497014 395818
rect 496394 395498 496426 395734
rect 496662 395498 496746 395734
rect 496982 395498 497014 395734
rect 496394 362054 497014 395498
rect 496394 361818 496426 362054
rect 496662 361818 496746 362054
rect 496982 361818 497014 362054
rect 496394 361734 497014 361818
rect 496394 361498 496426 361734
rect 496662 361498 496746 361734
rect 496982 361498 497014 361734
rect 496394 328054 497014 361498
rect 496394 327818 496426 328054
rect 496662 327818 496746 328054
rect 496982 327818 497014 328054
rect 496394 327734 497014 327818
rect 496394 327498 496426 327734
rect 496662 327498 496746 327734
rect 496982 327498 497014 327734
rect 496394 294054 497014 327498
rect 496394 293818 496426 294054
rect 496662 293818 496746 294054
rect 496982 293818 497014 294054
rect 496394 293734 497014 293818
rect 496394 293498 496426 293734
rect 496662 293498 496746 293734
rect 496982 293498 497014 293734
rect 496394 260054 497014 293498
rect 496394 259818 496426 260054
rect 496662 259818 496746 260054
rect 496982 259818 497014 260054
rect 496394 259734 497014 259818
rect 496394 259498 496426 259734
rect 496662 259498 496746 259734
rect 496982 259498 497014 259734
rect 496394 226054 497014 259498
rect 496394 225818 496426 226054
rect 496662 225818 496746 226054
rect 496982 225818 497014 226054
rect 496394 225734 497014 225818
rect 496394 225498 496426 225734
rect 496662 225498 496746 225734
rect 496982 225498 497014 225734
rect 496394 192054 497014 225498
rect 496394 191818 496426 192054
rect 496662 191818 496746 192054
rect 496982 191818 497014 192054
rect 496394 191734 497014 191818
rect 496394 191498 496426 191734
rect 496662 191498 496746 191734
rect 496982 191498 497014 191734
rect 496394 158054 497014 191498
rect 496394 157818 496426 158054
rect 496662 157818 496746 158054
rect 496982 157818 497014 158054
rect 496394 157734 497014 157818
rect 496394 157498 496426 157734
rect 496662 157498 496746 157734
rect 496982 157498 497014 157734
rect 496394 124054 497014 157498
rect 496394 123818 496426 124054
rect 496662 123818 496746 124054
rect 496982 123818 497014 124054
rect 496394 123734 497014 123818
rect 496394 123498 496426 123734
rect 496662 123498 496746 123734
rect 496982 123498 497014 123734
rect 496394 90054 497014 123498
rect 496394 89818 496426 90054
rect 496662 89818 496746 90054
rect 496982 89818 497014 90054
rect 496394 89734 497014 89818
rect 496394 89498 496426 89734
rect 496662 89498 496746 89734
rect 496982 89498 497014 89734
rect 496394 56054 497014 89498
rect 496394 55818 496426 56054
rect 496662 55818 496746 56054
rect 496982 55818 497014 56054
rect 496394 55734 497014 55818
rect 496394 55498 496426 55734
rect 496662 55498 496746 55734
rect 496982 55498 497014 55734
rect 496394 22054 497014 55498
rect 496394 21818 496426 22054
rect 496662 21818 496746 22054
rect 496982 21818 497014 22054
rect 496394 21734 497014 21818
rect 496394 21498 496426 21734
rect 496662 21498 496746 21734
rect 496982 21498 497014 21734
rect 496394 -5146 497014 21498
rect 496394 -5382 496426 -5146
rect 496662 -5382 496746 -5146
rect 496982 -5382 497014 -5146
rect 496394 -5466 497014 -5382
rect 496394 -5702 496426 -5466
rect 496662 -5702 496746 -5466
rect 496982 -5702 497014 -5466
rect 496394 -7654 497014 -5702
rect 500114 710598 500734 711590
rect 500114 710362 500146 710598
rect 500382 710362 500466 710598
rect 500702 710362 500734 710598
rect 500114 710278 500734 710362
rect 500114 710042 500146 710278
rect 500382 710042 500466 710278
rect 500702 710042 500734 710278
rect 500114 671774 500734 710042
rect 500114 671538 500146 671774
rect 500382 671538 500466 671774
rect 500702 671538 500734 671774
rect 500114 671454 500734 671538
rect 500114 671218 500146 671454
rect 500382 671218 500466 671454
rect 500702 671218 500734 671454
rect 500114 637774 500734 671218
rect 500114 637538 500146 637774
rect 500382 637538 500466 637774
rect 500702 637538 500734 637774
rect 500114 637454 500734 637538
rect 500114 637218 500146 637454
rect 500382 637218 500466 637454
rect 500702 637218 500734 637454
rect 500114 603774 500734 637218
rect 500114 603538 500146 603774
rect 500382 603538 500466 603774
rect 500702 603538 500734 603774
rect 500114 603454 500734 603538
rect 500114 603218 500146 603454
rect 500382 603218 500466 603454
rect 500702 603218 500734 603454
rect 500114 569774 500734 603218
rect 500114 569538 500146 569774
rect 500382 569538 500466 569774
rect 500702 569538 500734 569774
rect 500114 569454 500734 569538
rect 500114 569218 500146 569454
rect 500382 569218 500466 569454
rect 500702 569218 500734 569454
rect 500114 535774 500734 569218
rect 500114 535538 500146 535774
rect 500382 535538 500466 535774
rect 500702 535538 500734 535774
rect 500114 535454 500734 535538
rect 500114 535218 500146 535454
rect 500382 535218 500466 535454
rect 500702 535218 500734 535454
rect 500114 501774 500734 535218
rect 500114 501538 500146 501774
rect 500382 501538 500466 501774
rect 500702 501538 500734 501774
rect 500114 501454 500734 501538
rect 500114 501218 500146 501454
rect 500382 501218 500466 501454
rect 500702 501218 500734 501454
rect 500114 467774 500734 501218
rect 500114 467538 500146 467774
rect 500382 467538 500466 467774
rect 500702 467538 500734 467774
rect 500114 467454 500734 467538
rect 500114 467218 500146 467454
rect 500382 467218 500466 467454
rect 500702 467218 500734 467454
rect 500114 433774 500734 467218
rect 500114 433538 500146 433774
rect 500382 433538 500466 433774
rect 500702 433538 500734 433774
rect 500114 433454 500734 433538
rect 500114 433218 500146 433454
rect 500382 433218 500466 433454
rect 500702 433218 500734 433454
rect 500114 399774 500734 433218
rect 500114 399538 500146 399774
rect 500382 399538 500466 399774
rect 500702 399538 500734 399774
rect 500114 399454 500734 399538
rect 500114 399218 500146 399454
rect 500382 399218 500466 399454
rect 500702 399218 500734 399454
rect 500114 365774 500734 399218
rect 500114 365538 500146 365774
rect 500382 365538 500466 365774
rect 500702 365538 500734 365774
rect 500114 365454 500734 365538
rect 500114 365218 500146 365454
rect 500382 365218 500466 365454
rect 500702 365218 500734 365454
rect 500114 331774 500734 365218
rect 500114 331538 500146 331774
rect 500382 331538 500466 331774
rect 500702 331538 500734 331774
rect 500114 331454 500734 331538
rect 500114 331218 500146 331454
rect 500382 331218 500466 331454
rect 500702 331218 500734 331454
rect 500114 297774 500734 331218
rect 500114 297538 500146 297774
rect 500382 297538 500466 297774
rect 500702 297538 500734 297774
rect 500114 297454 500734 297538
rect 500114 297218 500146 297454
rect 500382 297218 500466 297454
rect 500702 297218 500734 297454
rect 500114 263774 500734 297218
rect 500114 263538 500146 263774
rect 500382 263538 500466 263774
rect 500702 263538 500734 263774
rect 500114 263454 500734 263538
rect 500114 263218 500146 263454
rect 500382 263218 500466 263454
rect 500702 263218 500734 263454
rect 500114 229774 500734 263218
rect 500114 229538 500146 229774
rect 500382 229538 500466 229774
rect 500702 229538 500734 229774
rect 500114 229454 500734 229538
rect 500114 229218 500146 229454
rect 500382 229218 500466 229454
rect 500702 229218 500734 229454
rect 500114 195774 500734 229218
rect 500114 195538 500146 195774
rect 500382 195538 500466 195774
rect 500702 195538 500734 195774
rect 500114 195454 500734 195538
rect 500114 195218 500146 195454
rect 500382 195218 500466 195454
rect 500702 195218 500734 195454
rect 500114 161774 500734 195218
rect 500114 161538 500146 161774
rect 500382 161538 500466 161774
rect 500702 161538 500734 161774
rect 500114 161454 500734 161538
rect 500114 161218 500146 161454
rect 500382 161218 500466 161454
rect 500702 161218 500734 161454
rect 500114 127774 500734 161218
rect 500114 127538 500146 127774
rect 500382 127538 500466 127774
rect 500702 127538 500734 127774
rect 500114 127454 500734 127538
rect 500114 127218 500146 127454
rect 500382 127218 500466 127454
rect 500702 127218 500734 127454
rect 500114 93774 500734 127218
rect 500114 93538 500146 93774
rect 500382 93538 500466 93774
rect 500702 93538 500734 93774
rect 500114 93454 500734 93538
rect 500114 93218 500146 93454
rect 500382 93218 500466 93454
rect 500702 93218 500734 93454
rect 500114 59774 500734 93218
rect 500114 59538 500146 59774
rect 500382 59538 500466 59774
rect 500702 59538 500734 59774
rect 500114 59454 500734 59538
rect 500114 59218 500146 59454
rect 500382 59218 500466 59454
rect 500702 59218 500734 59454
rect 500114 25774 500734 59218
rect 500114 25538 500146 25774
rect 500382 25538 500466 25774
rect 500702 25538 500734 25774
rect 500114 25454 500734 25538
rect 500114 25218 500146 25454
rect 500382 25218 500466 25454
rect 500702 25218 500734 25454
rect 500114 -6106 500734 25218
rect 500114 -6342 500146 -6106
rect 500382 -6342 500466 -6106
rect 500702 -6342 500734 -6106
rect 500114 -6426 500734 -6342
rect 500114 -6662 500146 -6426
rect 500382 -6662 500466 -6426
rect 500702 -6662 500734 -6426
rect 500114 -7654 500734 -6662
rect 503834 711558 504454 711590
rect 503834 711322 503866 711558
rect 504102 711322 504186 711558
rect 504422 711322 504454 711558
rect 503834 711238 504454 711322
rect 503834 711002 503866 711238
rect 504102 711002 504186 711238
rect 504422 711002 504454 711238
rect 503834 675494 504454 711002
rect 503834 675258 503866 675494
rect 504102 675258 504186 675494
rect 504422 675258 504454 675494
rect 503834 675174 504454 675258
rect 503834 674938 503866 675174
rect 504102 674938 504186 675174
rect 504422 674938 504454 675174
rect 503834 641494 504454 674938
rect 503834 641258 503866 641494
rect 504102 641258 504186 641494
rect 504422 641258 504454 641494
rect 503834 641174 504454 641258
rect 503834 640938 503866 641174
rect 504102 640938 504186 641174
rect 504422 640938 504454 641174
rect 503834 607494 504454 640938
rect 503834 607258 503866 607494
rect 504102 607258 504186 607494
rect 504422 607258 504454 607494
rect 503834 607174 504454 607258
rect 503834 606938 503866 607174
rect 504102 606938 504186 607174
rect 504422 606938 504454 607174
rect 503834 573494 504454 606938
rect 503834 573258 503866 573494
rect 504102 573258 504186 573494
rect 504422 573258 504454 573494
rect 503834 573174 504454 573258
rect 503834 572938 503866 573174
rect 504102 572938 504186 573174
rect 504422 572938 504454 573174
rect 503834 539494 504454 572938
rect 503834 539258 503866 539494
rect 504102 539258 504186 539494
rect 504422 539258 504454 539494
rect 503834 539174 504454 539258
rect 503834 538938 503866 539174
rect 504102 538938 504186 539174
rect 504422 538938 504454 539174
rect 503834 505494 504454 538938
rect 503834 505258 503866 505494
rect 504102 505258 504186 505494
rect 504422 505258 504454 505494
rect 503834 505174 504454 505258
rect 503834 504938 503866 505174
rect 504102 504938 504186 505174
rect 504422 504938 504454 505174
rect 503834 471494 504454 504938
rect 503834 471258 503866 471494
rect 504102 471258 504186 471494
rect 504422 471258 504454 471494
rect 503834 471174 504454 471258
rect 503834 470938 503866 471174
rect 504102 470938 504186 471174
rect 504422 470938 504454 471174
rect 503834 437494 504454 470938
rect 503834 437258 503866 437494
rect 504102 437258 504186 437494
rect 504422 437258 504454 437494
rect 503834 437174 504454 437258
rect 503834 436938 503866 437174
rect 504102 436938 504186 437174
rect 504422 436938 504454 437174
rect 503834 403494 504454 436938
rect 503834 403258 503866 403494
rect 504102 403258 504186 403494
rect 504422 403258 504454 403494
rect 503834 403174 504454 403258
rect 503834 402938 503866 403174
rect 504102 402938 504186 403174
rect 504422 402938 504454 403174
rect 503834 369494 504454 402938
rect 503834 369258 503866 369494
rect 504102 369258 504186 369494
rect 504422 369258 504454 369494
rect 503834 369174 504454 369258
rect 503834 368938 503866 369174
rect 504102 368938 504186 369174
rect 504422 368938 504454 369174
rect 503834 335494 504454 368938
rect 503834 335258 503866 335494
rect 504102 335258 504186 335494
rect 504422 335258 504454 335494
rect 503834 335174 504454 335258
rect 503834 334938 503866 335174
rect 504102 334938 504186 335174
rect 504422 334938 504454 335174
rect 503834 301494 504454 334938
rect 503834 301258 503866 301494
rect 504102 301258 504186 301494
rect 504422 301258 504454 301494
rect 503834 301174 504454 301258
rect 503834 300938 503866 301174
rect 504102 300938 504186 301174
rect 504422 300938 504454 301174
rect 503834 267494 504454 300938
rect 503834 267258 503866 267494
rect 504102 267258 504186 267494
rect 504422 267258 504454 267494
rect 503834 267174 504454 267258
rect 503834 266938 503866 267174
rect 504102 266938 504186 267174
rect 504422 266938 504454 267174
rect 503834 233494 504454 266938
rect 503834 233258 503866 233494
rect 504102 233258 504186 233494
rect 504422 233258 504454 233494
rect 503834 233174 504454 233258
rect 503834 232938 503866 233174
rect 504102 232938 504186 233174
rect 504422 232938 504454 233174
rect 503834 199494 504454 232938
rect 503834 199258 503866 199494
rect 504102 199258 504186 199494
rect 504422 199258 504454 199494
rect 503834 199174 504454 199258
rect 503834 198938 503866 199174
rect 504102 198938 504186 199174
rect 504422 198938 504454 199174
rect 503834 165494 504454 198938
rect 503834 165258 503866 165494
rect 504102 165258 504186 165494
rect 504422 165258 504454 165494
rect 503834 165174 504454 165258
rect 503834 164938 503866 165174
rect 504102 164938 504186 165174
rect 504422 164938 504454 165174
rect 503834 131494 504454 164938
rect 503834 131258 503866 131494
rect 504102 131258 504186 131494
rect 504422 131258 504454 131494
rect 503834 131174 504454 131258
rect 503834 130938 503866 131174
rect 504102 130938 504186 131174
rect 504422 130938 504454 131174
rect 503834 97494 504454 130938
rect 503834 97258 503866 97494
rect 504102 97258 504186 97494
rect 504422 97258 504454 97494
rect 503834 97174 504454 97258
rect 503834 96938 503866 97174
rect 504102 96938 504186 97174
rect 504422 96938 504454 97174
rect 503834 63494 504454 96938
rect 503834 63258 503866 63494
rect 504102 63258 504186 63494
rect 504422 63258 504454 63494
rect 503834 63174 504454 63258
rect 503834 62938 503866 63174
rect 504102 62938 504186 63174
rect 504422 62938 504454 63174
rect 503834 29494 504454 62938
rect 503834 29258 503866 29494
rect 504102 29258 504186 29494
rect 504422 29258 504454 29494
rect 503834 29174 504454 29258
rect 503834 28938 503866 29174
rect 504102 28938 504186 29174
rect 504422 28938 504454 29174
rect 503834 -7066 504454 28938
rect 503834 -7302 503866 -7066
rect 504102 -7302 504186 -7066
rect 504422 -7302 504454 -7066
rect 503834 -7386 504454 -7302
rect 503834 -7622 503866 -7386
rect 504102 -7622 504186 -7386
rect 504422 -7622 504454 -7386
rect 503834 -7654 504454 -7622
rect 511794 704838 512414 711590
rect 511794 704602 511826 704838
rect 512062 704602 512146 704838
rect 512382 704602 512414 704838
rect 511794 704518 512414 704602
rect 511794 704282 511826 704518
rect 512062 704282 512146 704518
rect 512382 704282 512414 704518
rect 511794 683454 512414 704282
rect 511794 683218 511826 683454
rect 512062 683218 512146 683454
rect 512382 683218 512414 683454
rect 511794 683134 512414 683218
rect 511794 682898 511826 683134
rect 512062 682898 512146 683134
rect 512382 682898 512414 683134
rect 511794 649454 512414 682898
rect 511794 649218 511826 649454
rect 512062 649218 512146 649454
rect 512382 649218 512414 649454
rect 511794 649134 512414 649218
rect 511794 648898 511826 649134
rect 512062 648898 512146 649134
rect 512382 648898 512414 649134
rect 511794 615454 512414 648898
rect 511794 615218 511826 615454
rect 512062 615218 512146 615454
rect 512382 615218 512414 615454
rect 511794 615134 512414 615218
rect 511794 614898 511826 615134
rect 512062 614898 512146 615134
rect 512382 614898 512414 615134
rect 511794 581454 512414 614898
rect 511794 581218 511826 581454
rect 512062 581218 512146 581454
rect 512382 581218 512414 581454
rect 511794 581134 512414 581218
rect 511794 580898 511826 581134
rect 512062 580898 512146 581134
rect 512382 580898 512414 581134
rect 511794 547454 512414 580898
rect 511794 547218 511826 547454
rect 512062 547218 512146 547454
rect 512382 547218 512414 547454
rect 511794 547134 512414 547218
rect 511794 546898 511826 547134
rect 512062 546898 512146 547134
rect 512382 546898 512414 547134
rect 511794 513454 512414 546898
rect 511794 513218 511826 513454
rect 512062 513218 512146 513454
rect 512382 513218 512414 513454
rect 511794 513134 512414 513218
rect 511794 512898 511826 513134
rect 512062 512898 512146 513134
rect 512382 512898 512414 513134
rect 511794 479454 512414 512898
rect 511794 479218 511826 479454
rect 512062 479218 512146 479454
rect 512382 479218 512414 479454
rect 511794 479134 512414 479218
rect 511794 478898 511826 479134
rect 512062 478898 512146 479134
rect 512382 478898 512414 479134
rect 511794 445454 512414 478898
rect 511794 445218 511826 445454
rect 512062 445218 512146 445454
rect 512382 445218 512414 445454
rect 511794 445134 512414 445218
rect 511794 444898 511826 445134
rect 512062 444898 512146 445134
rect 512382 444898 512414 445134
rect 511794 411454 512414 444898
rect 511794 411218 511826 411454
rect 512062 411218 512146 411454
rect 512382 411218 512414 411454
rect 511794 411134 512414 411218
rect 511794 410898 511826 411134
rect 512062 410898 512146 411134
rect 512382 410898 512414 411134
rect 511794 377454 512414 410898
rect 511794 377218 511826 377454
rect 512062 377218 512146 377454
rect 512382 377218 512414 377454
rect 511794 377134 512414 377218
rect 511794 376898 511826 377134
rect 512062 376898 512146 377134
rect 512382 376898 512414 377134
rect 511794 343454 512414 376898
rect 511794 343218 511826 343454
rect 512062 343218 512146 343454
rect 512382 343218 512414 343454
rect 511794 343134 512414 343218
rect 511794 342898 511826 343134
rect 512062 342898 512146 343134
rect 512382 342898 512414 343134
rect 511794 309454 512414 342898
rect 511794 309218 511826 309454
rect 512062 309218 512146 309454
rect 512382 309218 512414 309454
rect 511794 309134 512414 309218
rect 511794 308898 511826 309134
rect 512062 308898 512146 309134
rect 512382 308898 512414 309134
rect 511794 275454 512414 308898
rect 511794 275218 511826 275454
rect 512062 275218 512146 275454
rect 512382 275218 512414 275454
rect 511794 275134 512414 275218
rect 511794 274898 511826 275134
rect 512062 274898 512146 275134
rect 512382 274898 512414 275134
rect 511794 241454 512414 274898
rect 511794 241218 511826 241454
rect 512062 241218 512146 241454
rect 512382 241218 512414 241454
rect 511794 241134 512414 241218
rect 511794 240898 511826 241134
rect 512062 240898 512146 241134
rect 512382 240898 512414 241134
rect 511794 207454 512414 240898
rect 511794 207218 511826 207454
rect 512062 207218 512146 207454
rect 512382 207218 512414 207454
rect 511794 207134 512414 207218
rect 511794 206898 511826 207134
rect 512062 206898 512146 207134
rect 512382 206898 512414 207134
rect 511794 173454 512414 206898
rect 511794 173218 511826 173454
rect 512062 173218 512146 173454
rect 512382 173218 512414 173454
rect 511794 173134 512414 173218
rect 511794 172898 511826 173134
rect 512062 172898 512146 173134
rect 512382 172898 512414 173134
rect 511794 139454 512414 172898
rect 511794 139218 511826 139454
rect 512062 139218 512146 139454
rect 512382 139218 512414 139454
rect 511794 139134 512414 139218
rect 511794 138898 511826 139134
rect 512062 138898 512146 139134
rect 512382 138898 512414 139134
rect 511794 105454 512414 138898
rect 511794 105218 511826 105454
rect 512062 105218 512146 105454
rect 512382 105218 512414 105454
rect 511794 105134 512414 105218
rect 511794 104898 511826 105134
rect 512062 104898 512146 105134
rect 512382 104898 512414 105134
rect 511794 71454 512414 104898
rect 511794 71218 511826 71454
rect 512062 71218 512146 71454
rect 512382 71218 512414 71454
rect 511794 71134 512414 71218
rect 511794 70898 511826 71134
rect 512062 70898 512146 71134
rect 512382 70898 512414 71134
rect 511794 37454 512414 70898
rect 511794 37218 511826 37454
rect 512062 37218 512146 37454
rect 512382 37218 512414 37454
rect 511794 37134 512414 37218
rect 511794 36898 511826 37134
rect 512062 36898 512146 37134
rect 512382 36898 512414 37134
rect 511794 3454 512414 36898
rect 511794 3218 511826 3454
rect 512062 3218 512146 3454
rect 512382 3218 512414 3454
rect 511794 3134 512414 3218
rect 511794 2898 511826 3134
rect 512062 2898 512146 3134
rect 512382 2898 512414 3134
rect 511794 -346 512414 2898
rect 511794 -582 511826 -346
rect 512062 -582 512146 -346
rect 512382 -582 512414 -346
rect 511794 -666 512414 -582
rect 511794 -902 511826 -666
rect 512062 -902 512146 -666
rect 512382 -902 512414 -666
rect 511794 -7654 512414 -902
rect 515514 705798 516134 711590
rect 515514 705562 515546 705798
rect 515782 705562 515866 705798
rect 516102 705562 516134 705798
rect 515514 705478 516134 705562
rect 515514 705242 515546 705478
rect 515782 705242 515866 705478
rect 516102 705242 516134 705478
rect 515514 687174 516134 705242
rect 515514 686938 515546 687174
rect 515782 686938 515866 687174
rect 516102 686938 516134 687174
rect 515514 686854 516134 686938
rect 515514 686618 515546 686854
rect 515782 686618 515866 686854
rect 516102 686618 516134 686854
rect 515514 653174 516134 686618
rect 515514 652938 515546 653174
rect 515782 652938 515866 653174
rect 516102 652938 516134 653174
rect 515514 652854 516134 652938
rect 515514 652618 515546 652854
rect 515782 652618 515866 652854
rect 516102 652618 516134 652854
rect 515514 619174 516134 652618
rect 515514 618938 515546 619174
rect 515782 618938 515866 619174
rect 516102 618938 516134 619174
rect 515514 618854 516134 618938
rect 515514 618618 515546 618854
rect 515782 618618 515866 618854
rect 516102 618618 516134 618854
rect 515514 585174 516134 618618
rect 515514 584938 515546 585174
rect 515782 584938 515866 585174
rect 516102 584938 516134 585174
rect 515514 584854 516134 584938
rect 515514 584618 515546 584854
rect 515782 584618 515866 584854
rect 516102 584618 516134 584854
rect 515514 551174 516134 584618
rect 515514 550938 515546 551174
rect 515782 550938 515866 551174
rect 516102 550938 516134 551174
rect 515514 550854 516134 550938
rect 515514 550618 515546 550854
rect 515782 550618 515866 550854
rect 516102 550618 516134 550854
rect 515514 517174 516134 550618
rect 515514 516938 515546 517174
rect 515782 516938 515866 517174
rect 516102 516938 516134 517174
rect 515514 516854 516134 516938
rect 515514 516618 515546 516854
rect 515782 516618 515866 516854
rect 516102 516618 516134 516854
rect 515514 483174 516134 516618
rect 515514 482938 515546 483174
rect 515782 482938 515866 483174
rect 516102 482938 516134 483174
rect 515514 482854 516134 482938
rect 515514 482618 515546 482854
rect 515782 482618 515866 482854
rect 516102 482618 516134 482854
rect 515514 449174 516134 482618
rect 515514 448938 515546 449174
rect 515782 448938 515866 449174
rect 516102 448938 516134 449174
rect 515514 448854 516134 448938
rect 515514 448618 515546 448854
rect 515782 448618 515866 448854
rect 516102 448618 516134 448854
rect 515514 415174 516134 448618
rect 515514 414938 515546 415174
rect 515782 414938 515866 415174
rect 516102 414938 516134 415174
rect 515514 414854 516134 414938
rect 515514 414618 515546 414854
rect 515782 414618 515866 414854
rect 516102 414618 516134 414854
rect 515514 381174 516134 414618
rect 515514 380938 515546 381174
rect 515782 380938 515866 381174
rect 516102 380938 516134 381174
rect 515514 380854 516134 380938
rect 515514 380618 515546 380854
rect 515782 380618 515866 380854
rect 516102 380618 516134 380854
rect 515514 347174 516134 380618
rect 515514 346938 515546 347174
rect 515782 346938 515866 347174
rect 516102 346938 516134 347174
rect 515514 346854 516134 346938
rect 515514 346618 515546 346854
rect 515782 346618 515866 346854
rect 516102 346618 516134 346854
rect 515514 313174 516134 346618
rect 515514 312938 515546 313174
rect 515782 312938 515866 313174
rect 516102 312938 516134 313174
rect 515514 312854 516134 312938
rect 515514 312618 515546 312854
rect 515782 312618 515866 312854
rect 516102 312618 516134 312854
rect 515514 279174 516134 312618
rect 515514 278938 515546 279174
rect 515782 278938 515866 279174
rect 516102 278938 516134 279174
rect 515514 278854 516134 278938
rect 515514 278618 515546 278854
rect 515782 278618 515866 278854
rect 516102 278618 516134 278854
rect 515514 245174 516134 278618
rect 515514 244938 515546 245174
rect 515782 244938 515866 245174
rect 516102 244938 516134 245174
rect 515514 244854 516134 244938
rect 515514 244618 515546 244854
rect 515782 244618 515866 244854
rect 516102 244618 516134 244854
rect 515514 211174 516134 244618
rect 515514 210938 515546 211174
rect 515782 210938 515866 211174
rect 516102 210938 516134 211174
rect 515514 210854 516134 210938
rect 515514 210618 515546 210854
rect 515782 210618 515866 210854
rect 516102 210618 516134 210854
rect 515514 177174 516134 210618
rect 515514 176938 515546 177174
rect 515782 176938 515866 177174
rect 516102 176938 516134 177174
rect 515514 176854 516134 176938
rect 515514 176618 515546 176854
rect 515782 176618 515866 176854
rect 516102 176618 516134 176854
rect 515514 143174 516134 176618
rect 515514 142938 515546 143174
rect 515782 142938 515866 143174
rect 516102 142938 516134 143174
rect 515514 142854 516134 142938
rect 515514 142618 515546 142854
rect 515782 142618 515866 142854
rect 516102 142618 516134 142854
rect 515514 109174 516134 142618
rect 515514 108938 515546 109174
rect 515782 108938 515866 109174
rect 516102 108938 516134 109174
rect 515514 108854 516134 108938
rect 515514 108618 515546 108854
rect 515782 108618 515866 108854
rect 516102 108618 516134 108854
rect 515514 75174 516134 108618
rect 515514 74938 515546 75174
rect 515782 74938 515866 75174
rect 516102 74938 516134 75174
rect 515514 74854 516134 74938
rect 515514 74618 515546 74854
rect 515782 74618 515866 74854
rect 516102 74618 516134 74854
rect 515514 41174 516134 74618
rect 515514 40938 515546 41174
rect 515782 40938 515866 41174
rect 516102 40938 516134 41174
rect 515514 40854 516134 40938
rect 515514 40618 515546 40854
rect 515782 40618 515866 40854
rect 516102 40618 516134 40854
rect 515514 7174 516134 40618
rect 515514 6938 515546 7174
rect 515782 6938 515866 7174
rect 516102 6938 516134 7174
rect 515514 6854 516134 6938
rect 515514 6618 515546 6854
rect 515782 6618 515866 6854
rect 516102 6618 516134 6854
rect 515514 -1306 516134 6618
rect 515514 -1542 515546 -1306
rect 515782 -1542 515866 -1306
rect 516102 -1542 516134 -1306
rect 515514 -1626 516134 -1542
rect 515514 -1862 515546 -1626
rect 515782 -1862 515866 -1626
rect 516102 -1862 516134 -1626
rect 515514 -7654 516134 -1862
rect 519234 706758 519854 711590
rect 519234 706522 519266 706758
rect 519502 706522 519586 706758
rect 519822 706522 519854 706758
rect 519234 706438 519854 706522
rect 519234 706202 519266 706438
rect 519502 706202 519586 706438
rect 519822 706202 519854 706438
rect 519234 690894 519854 706202
rect 519234 690658 519266 690894
rect 519502 690658 519586 690894
rect 519822 690658 519854 690894
rect 519234 690574 519854 690658
rect 519234 690338 519266 690574
rect 519502 690338 519586 690574
rect 519822 690338 519854 690574
rect 519234 656894 519854 690338
rect 519234 656658 519266 656894
rect 519502 656658 519586 656894
rect 519822 656658 519854 656894
rect 519234 656574 519854 656658
rect 519234 656338 519266 656574
rect 519502 656338 519586 656574
rect 519822 656338 519854 656574
rect 519234 622894 519854 656338
rect 519234 622658 519266 622894
rect 519502 622658 519586 622894
rect 519822 622658 519854 622894
rect 519234 622574 519854 622658
rect 519234 622338 519266 622574
rect 519502 622338 519586 622574
rect 519822 622338 519854 622574
rect 519234 588894 519854 622338
rect 519234 588658 519266 588894
rect 519502 588658 519586 588894
rect 519822 588658 519854 588894
rect 519234 588574 519854 588658
rect 519234 588338 519266 588574
rect 519502 588338 519586 588574
rect 519822 588338 519854 588574
rect 519234 554894 519854 588338
rect 519234 554658 519266 554894
rect 519502 554658 519586 554894
rect 519822 554658 519854 554894
rect 519234 554574 519854 554658
rect 519234 554338 519266 554574
rect 519502 554338 519586 554574
rect 519822 554338 519854 554574
rect 519234 520894 519854 554338
rect 519234 520658 519266 520894
rect 519502 520658 519586 520894
rect 519822 520658 519854 520894
rect 519234 520574 519854 520658
rect 519234 520338 519266 520574
rect 519502 520338 519586 520574
rect 519822 520338 519854 520574
rect 519234 486894 519854 520338
rect 519234 486658 519266 486894
rect 519502 486658 519586 486894
rect 519822 486658 519854 486894
rect 519234 486574 519854 486658
rect 519234 486338 519266 486574
rect 519502 486338 519586 486574
rect 519822 486338 519854 486574
rect 519234 452894 519854 486338
rect 519234 452658 519266 452894
rect 519502 452658 519586 452894
rect 519822 452658 519854 452894
rect 519234 452574 519854 452658
rect 519234 452338 519266 452574
rect 519502 452338 519586 452574
rect 519822 452338 519854 452574
rect 519234 418894 519854 452338
rect 519234 418658 519266 418894
rect 519502 418658 519586 418894
rect 519822 418658 519854 418894
rect 519234 418574 519854 418658
rect 519234 418338 519266 418574
rect 519502 418338 519586 418574
rect 519822 418338 519854 418574
rect 519234 384894 519854 418338
rect 519234 384658 519266 384894
rect 519502 384658 519586 384894
rect 519822 384658 519854 384894
rect 519234 384574 519854 384658
rect 519234 384338 519266 384574
rect 519502 384338 519586 384574
rect 519822 384338 519854 384574
rect 519234 350894 519854 384338
rect 519234 350658 519266 350894
rect 519502 350658 519586 350894
rect 519822 350658 519854 350894
rect 519234 350574 519854 350658
rect 519234 350338 519266 350574
rect 519502 350338 519586 350574
rect 519822 350338 519854 350574
rect 519234 316894 519854 350338
rect 519234 316658 519266 316894
rect 519502 316658 519586 316894
rect 519822 316658 519854 316894
rect 519234 316574 519854 316658
rect 519234 316338 519266 316574
rect 519502 316338 519586 316574
rect 519822 316338 519854 316574
rect 519234 282894 519854 316338
rect 519234 282658 519266 282894
rect 519502 282658 519586 282894
rect 519822 282658 519854 282894
rect 519234 282574 519854 282658
rect 519234 282338 519266 282574
rect 519502 282338 519586 282574
rect 519822 282338 519854 282574
rect 519234 248894 519854 282338
rect 519234 248658 519266 248894
rect 519502 248658 519586 248894
rect 519822 248658 519854 248894
rect 519234 248574 519854 248658
rect 519234 248338 519266 248574
rect 519502 248338 519586 248574
rect 519822 248338 519854 248574
rect 519234 214894 519854 248338
rect 519234 214658 519266 214894
rect 519502 214658 519586 214894
rect 519822 214658 519854 214894
rect 519234 214574 519854 214658
rect 519234 214338 519266 214574
rect 519502 214338 519586 214574
rect 519822 214338 519854 214574
rect 519234 180894 519854 214338
rect 519234 180658 519266 180894
rect 519502 180658 519586 180894
rect 519822 180658 519854 180894
rect 519234 180574 519854 180658
rect 519234 180338 519266 180574
rect 519502 180338 519586 180574
rect 519822 180338 519854 180574
rect 519234 146894 519854 180338
rect 519234 146658 519266 146894
rect 519502 146658 519586 146894
rect 519822 146658 519854 146894
rect 519234 146574 519854 146658
rect 519234 146338 519266 146574
rect 519502 146338 519586 146574
rect 519822 146338 519854 146574
rect 519234 112894 519854 146338
rect 519234 112658 519266 112894
rect 519502 112658 519586 112894
rect 519822 112658 519854 112894
rect 519234 112574 519854 112658
rect 519234 112338 519266 112574
rect 519502 112338 519586 112574
rect 519822 112338 519854 112574
rect 519234 78894 519854 112338
rect 519234 78658 519266 78894
rect 519502 78658 519586 78894
rect 519822 78658 519854 78894
rect 519234 78574 519854 78658
rect 519234 78338 519266 78574
rect 519502 78338 519586 78574
rect 519822 78338 519854 78574
rect 519234 44894 519854 78338
rect 519234 44658 519266 44894
rect 519502 44658 519586 44894
rect 519822 44658 519854 44894
rect 519234 44574 519854 44658
rect 519234 44338 519266 44574
rect 519502 44338 519586 44574
rect 519822 44338 519854 44574
rect 519234 10894 519854 44338
rect 519234 10658 519266 10894
rect 519502 10658 519586 10894
rect 519822 10658 519854 10894
rect 519234 10574 519854 10658
rect 519234 10338 519266 10574
rect 519502 10338 519586 10574
rect 519822 10338 519854 10574
rect 519234 -2266 519854 10338
rect 519234 -2502 519266 -2266
rect 519502 -2502 519586 -2266
rect 519822 -2502 519854 -2266
rect 519234 -2586 519854 -2502
rect 519234 -2822 519266 -2586
rect 519502 -2822 519586 -2586
rect 519822 -2822 519854 -2586
rect 519234 -7654 519854 -2822
rect 522954 707718 523574 711590
rect 522954 707482 522986 707718
rect 523222 707482 523306 707718
rect 523542 707482 523574 707718
rect 522954 707398 523574 707482
rect 522954 707162 522986 707398
rect 523222 707162 523306 707398
rect 523542 707162 523574 707398
rect 522954 694614 523574 707162
rect 522954 694378 522986 694614
rect 523222 694378 523306 694614
rect 523542 694378 523574 694614
rect 522954 694294 523574 694378
rect 522954 694058 522986 694294
rect 523222 694058 523306 694294
rect 523542 694058 523574 694294
rect 522954 660614 523574 694058
rect 522954 660378 522986 660614
rect 523222 660378 523306 660614
rect 523542 660378 523574 660614
rect 522954 660294 523574 660378
rect 522954 660058 522986 660294
rect 523222 660058 523306 660294
rect 523542 660058 523574 660294
rect 522954 626614 523574 660058
rect 522954 626378 522986 626614
rect 523222 626378 523306 626614
rect 523542 626378 523574 626614
rect 522954 626294 523574 626378
rect 522954 626058 522986 626294
rect 523222 626058 523306 626294
rect 523542 626058 523574 626294
rect 522954 592614 523574 626058
rect 522954 592378 522986 592614
rect 523222 592378 523306 592614
rect 523542 592378 523574 592614
rect 522954 592294 523574 592378
rect 522954 592058 522986 592294
rect 523222 592058 523306 592294
rect 523542 592058 523574 592294
rect 522954 558614 523574 592058
rect 522954 558378 522986 558614
rect 523222 558378 523306 558614
rect 523542 558378 523574 558614
rect 522954 558294 523574 558378
rect 522954 558058 522986 558294
rect 523222 558058 523306 558294
rect 523542 558058 523574 558294
rect 522954 524614 523574 558058
rect 522954 524378 522986 524614
rect 523222 524378 523306 524614
rect 523542 524378 523574 524614
rect 522954 524294 523574 524378
rect 522954 524058 522986 524294
rect 523222 524058 523306 524294
rect 523542 524058 523574 524294
rect 522954 490614 523574 524058
rect 522954 490378 522986 490614
rect 523222 490378 523306 490614
rect 523542 490378 523574 490614
rect 522954 490294 523574 490378
rect 522954 490058 522986 490294
rect 523222 490058 523306 490294
rect 523542 490058 523574 490294
rect 522954 456614 523574 490058
rect 522954 456378 522986 456614
rect 523222 456378 523306 456614
rect 523542 456378 523574 456614
rect 522954 456294 523574 456378
rect 522954 456058 522986 456294
rect 523222 456058 523306 456294
rect 523542 456058 523574 456294
rect 522954 422614 523574 456058
rect 522954 422378 522986 422614
rect 523222 422378 523306 422614
rect 523542 422378 523574 422614
rect 522954 422294 523574 422378
rect 522954 422058 522986 422294
rect 523222 422058 523306 422294
rect 523542 422058 523574 422294
rect 522954 388614 523574 422058
rect 522954 388378 522986 388614
rect 523222 388378 523306 388614
rect 523542 388378 523574 388614
rect 522954 388294 523574 388378
rect 522954 388058 522986 388294
rect 523222 388058 523306 388294
rect 523542 388058 523574 388294
rect 522954 354614 523574 388058
rect 522954 354378 522986 354614
rect 523222 354378 523306 354614
rect 523542 354378 523574 354614
rect 522954 354294 523574 354378
rect 522954 354058 522986 354294
rect 523222 354058 523306 354294
rect 523542 354058 523574 354294
rect 522954 320614 523574 354058
rect 522954 320378 522986 320614
rect 523222 320378 523306 320614
rect 523542 320378 523574 320614
rect 522954 320294 523574 320378
rect 522954 320058 522986 320294
rect 523222 320058 523306 320294
rect 523542 320058 523574 320294
rect 522954 286614 523574 320058
rect 522954 286378 522986 286614
rect 523222 286378 523306 286614
rect 523542 286378 523574 286614
rect 522954 286294 523574 286378
rect 522954 286058 522986 286294
rect 523222 286058 523306 286294
rect 523542 286058 523574 286294
rect 522954 252614 523574 286058
rect 522954 252378 522986 252614
rect 523222 252378 523306 252614
rect 523542 252378 523574 252614
rect 522954 252294 523574 252378
rect 522954 252058 522986 252294
rect 523222 252058 523306 252294
rect 523542 252058 523574 252294
rect 522954 218614 523574 252058
rect 522954 218378 522986 218614
rect 523222 218378 523306 218614
rect 523542 218378 523574 218614
rect 522954 218294 523574 218378
rect 522954 218058 522986 218294
rect 523222 218058 523306 218294
rect 523542 218058 523574 218294
rect 522954 184614 523574 218058
rect 522954 184378 522986 184614
rect 523222 184378 523306 184614
rect 523542 184378 523574 184614
rect 522954 184294 523574 184378
rect 522954 184058 522986 184294
rect 523222 184058 523306 184294
rect 523542 184058 523574 184294
rect 522954 150614 523574 184058
rect 522954 150378 522986 150614
rect 523222 150378 523306 150614
rect 523542 150378 523574 150614
rect 522954 150294 523574 150378
rect 522954 150058 522986 150294
rect 523222 150058 523306 150294
rect 523542 150058 523574 150294
rect 522954 116614 523574 150058
rect 522954 116378 522986 116614
rect 523222 116378 523306 116614
rect 523542 116378 523574 116614
rect 522954 116294 523574 116378
rect 522954 116058 522986 116294
rect 523222 116058 523306 116294
rect 523542 116058 523574 116294
rect 522954 82614 523574 116058
rect 522954 82378 522986 82614
rect 523222 82378 523306 82614
rect 523542 82378 523574 82614
rect 522954 82294 523574 82378
rect 522954 82058 522986 82294
rect 523222 82058 523306 82294
rect 523542 82058 523574 82294
rect 522954 48614 523574 82058
rect 522954 48378 522986 48614
rect 523222 48378 523306 48614
rect 523542 48378 523574 48614
rect 522954 48294 523574 48378
rect 522954 48058 522986 48294
rect 523222 48058 523306 48294
rect 523542 48058 523574 48294
rect 522954 14614 523574 48058
rect 522954 14378 522986 14614
rect 523222 14378 523306 14614
rect 523542 14378 523574 14614
rect 522954 14294 523574 14378
rect 522954 14058 522986 14294
rect 523222 14058 523306 14294
rect 523542 14058 523574 14294
rect 522954 -3226 523574 14058
rect 522954 -3462 522986 -3226
rect 523222 -3462 523306 -3226
rect 523542 -3462 523574 -3226
rect 522954 -3546 523574 -3462
rect 522954 -3782 522986 -3546
rect 523222 -3782 523306 -3546
rect 523542 -3782 523574 -3546
rect 522954 -7654 523574 -3782
rect 526674 708678 527294 711590
rect 526674 708442 526706 708678
rect 526942 708442 527026 708678
rect 527262 708442 527294 708678
rect 526674 708358 527294 708442
rect 526674 708122 526706 708358
rect 526942 708122 527026 708358
rect 527262 708122 527294 708358
rect 526674 698334 527294 708122
rect 526674 698098 526706 698334
rect 526942 698098 527026 698334
rect 527262 698098 527294 698334
rect 526674 698014 527294 698098
rect 526674 697778 526706 698014
rect 526942 697778 527026 698014
rect 527262 697778 527294 698014
rect 526674 664334 527294 697778
rect 526674 664098 526706 664334
rect 526942 664098 527026 664334
rect 527262 664098 527294 664334
rect 526674 664014 527294 664098
rect 526674 663778 526706 664014
rect 526942 663778 527026 664014
rect 527262 663778 527294 664014
rect 526674 630334 527294 663778
rect 526674 630098 526706 630334
rect 526942 630098 527026 630334
rect 527262 630098 527294 630334
rect 526674 630014 527294 630098
rect 526674 629778 526706 630014
rect 526942 629778 527026 630014
rect 527262 629778 527294 630014
rect 526674 596334 527294 629778
rect 526674 596098 526706 596334
rect 526942 596098 527026 596334
rect 527262 596098 527294 596334
rect 526674 596014 527294 596098
rect 526674 595778 526706 596014
rect 526942 595778 527026 596014
rect 527262 595778 527294 596014
rect 526674 562334 527294 595778
rect 526674 562098 526706 562334
rect 526942 562098 527026 562334
rect 527262 562098 527294 562334
rect 526674 562014 527294 562098
rect 526674 561778 526706 562014
rect 526942 561778 527026 562014
rect 527262 561778 527294 562014
rect 526674 528334 527294 561778
rect 526674 528098 526706 528334
rect 526942 528098 527026 528334
rect 527262 528098 527294 528334
rect 526674 528014 527294 528098
rect 526674 527778 526706 528014
rect 526942 527778 527026 528014
rect 527262 527778 527294 528014
rect 526674 494334 527294 527778
rect 526674 494098 526706 494334
rect 526942 494098 527026 494334
rect 527262 494098 527294 494334
rect 526674 494014 527294 494098
rect 526674 493778 526706 494014
rect 526942 493778 527026 494014
rect 527262 493778 527294 494014
rect 526674 460334 527294 493778
rect 526674 460098 526706 460334
rect 526942 460098 527026 460334
rect 527262 460098 527294 460334
rect 526674 460014 527294 460098
rect 526674 459778 526706 460014
rect 526942 459778 527026 460014
rect 527262 459778 527294 460014
rect 526674 426334 527294 459778
rect 526674 426098 526706 426334
rect 526942 426098 527026 426334
rect 527262 426098 527294 426334
rect 526674 426014 527294 426098
rect 526674 425778 526706 426014
rect 526942 425778 527026 426014
rect 527262 425778 527294 426014
rect 526674 392334 527294 425778
rect 526674 392098 526706 392334
rect 526942 392098 527026 392334
rect 527262 392098 527294 392334
rect 526674 392014 527294 392098
rect 526674 391778 526706 392014
rect 526942 391778 527026 392014
rect 527262 391778 527294 392014
rect 526674 358334 527294 391778
rect 526674 358098 526706 358334
rect 526942 358098 527026 358334
rect 527262 358098 527294 358334
rect 526674 358014 527294 358098
rect 526674 357778 526706 358014
rect 526942 357778 527026 358014
rect 527262 357778 527294 358014
rect 526674 324334 527294 357778
rect 526674 324098 526706 324334
rect 526942 324098 527026 324334
rect 527262 324098 527294 324334
rect 526674 324014 527294 324098
rect 526674 323778 526706 324014
rect 526942 323778 527026 324014
rect 527262 323778 527294 324014
rect 526674 290334 527294 323778
rect 526674 290098 526706 290334
rect 526942 290098 527026 290334
rect 527262 290098 527294 290334
rect 526674 290014 527294 290098
rect 526674 289778 526706 290014
rect 526942 289778 527026 290014
rect 527262 289778 527294 290014
rect 526674 256334 527294 289778
rect 526674 256098 526706 256334
rect 526942 256098 527026 256334
rect 527262 256098 527294 256334
rect 526674 256014 527294 256098
rect 526674 255778 526706 256014
rect 526942 255778 527026 256014
rect 527262 255778 527294 256014
rect 526674 222334 527294 255778
rect 526674 222098 526706 222334
rect 526942 222098 527026 222334
rect 527262 222098 527294 222334
rect 526674 222014 527294 222098
rect 526674 221778 526706 222014
rect 526942 221778 527026 222014
rect 527262 221778 527294 222014
rect 526674 188334 527294 221778
rect 526674 188098 526706 188334
rect 526942 188098 527026 188334
rect 527262 188098 527294 188334
rect 526674 188014 527294 188098
rect 526674 187778 526706 188014
rect 526942 187778 527026 188014
rect 527262 187778 527294 188014
rect 526674 154334 527294 187778
rect 526674 154098 526706 154334
rect 526942 154098 527026 154334
rect 527262 154098 527294 154334
rect 526674 154014 527294 154098
rect 526674 153778 526706 154014
rect 526942 153778 527026 154014
rect 527262 153778 527294 154014
rect 526674 120334 527294 153778
rect 526674 120098 526706 120334
rect 526942 120098 527026 120334
rect 527262 120098 527294 120334
rect 526674 120014 527294 120098
rect 526674 119778 526706 120014
rect 526942 119778 527026 120014
rect 527262 119778 527294 120014
rect 526674 86334 527294 119778
rect 526674 86098 526706 86334
rect 526942 86098 527026 86334
rect 527262 86098 527294 86334
rect 526674 86014 527294 86098
rect 526674 85778 526706 86014
rect 526942 85778 527026 86014
rect 527262 85778 527294 86014
rect 526674 52334 527294 85778
rect 526674 52098 526706 52334
rect 526942 52098 527026 52334
rect 527262 52098 527294 52334
rect 526674 52014 527294 52098
rect 526674 51778 526706 52014
rect 526942 51778 527026 52014
rect 527262 51778 527294 52014
rect 526674 18334 527294 51778
rect 526674 18098 526706 18334
rect 526942 18098 527026 18334
rect 527262 18098 527294 18334
rect 526674 18014 527294 18098
rect 526674 17778 526706 18014
rect 526942 17778 527026 18014
rect 527262 17778 527294 18014
rect 526674 -4186 527294 17778
rect 526674 -4422 526706 -4186
rect 526942 -4422 527026 -4186
rect 527262 -4422 527294 -4186
rect 526674 -4506 527294 -4422
rect 526674 -4742 526706 -4506
rect 526942 -4742 527026 -4506
rect 527262 -4742 527294 -4506
rect 526674 -7654 527294 -4742
rect 530394 709638 531014 711590
rect 530394 709402 530426 709638
rect 530662 709402 530746 709638
rect 530982 709402 531014 709638
rect 530394 709318 531014 709402
rect 530394 709082 530426 709318
rect 530662 709082 530746 709318
rect 530982 709082 531014 709318
rect 530394 668054 531014 709082
rect 530394 667818 530426 668054
rect 530662 667818 530746 668054
rect 530982 667818 531014 668054
rect 530394 667734 531014 667818
rect 530394 667498 530426 667734
rect 530662 667498 530746 667734
rect 530982 667498 531014 667734
rect 530394 634054 531014 667498
rect 530394 633818 530426 634054
rect 530662 633818 530746 634054
rect 530982 633818 531014 634054
rect 530394 633734 531014 633818
rect 530394 633498 530426 633734
rect 530662 633498 530746 633734
rect 530982 633498 531014 633734
rect 530394 600054 531014 633498
rect 530394 599818 530426 600054
rect 530662 599818 530746 600054
rect 530982 599818 531014 600054
rect 530394 599734 531014 599818
rect 530394 599498 530426 599734
rect 530662 599498 530746 599734
rect 530982 599498 531014 599734
rect 530394 566054 531014 599498
rect 530394 565818 530426 566054
rect 530662 565818 530746 566054
rect 530982 565818 531014 566054
rect 530394 565734 531014 565818
rect 530394 565498 530426 565734
rect 530662 565498 530746 565734
rect 530982 565498 531014 565734
rect 530394 532054 531014 565498
rect 530394 531818 530426 532054
rect 530662 531818 530746 532054
rect 530982 531818 531014 532054
rect 530394 531734 531014 531818
rect 530394 531498 530426 531734
rect 530662 531498 530746 531734
rect 530982 531498 531014 531734
rect 530394 498054 531014 531498
rect 530394 497818 530426 498054
rect 530662 497818 530746 498054
rect 530982 497818 531014 498054
rect 530394 497734 531014 497818
rect 530394 497498 530426 497734
rect 530662 497498 530746 497734
rect 530982 497498 531014 497734
rect 530394 464054 531014 497498
rect 530394 463818 530426 464054
rect 530662 463818 530746 464054
rect 530982 463818 531014 464054
rect 530394 463734 531014 463818
rect 530394 463498 530426 463734
rect 530662 463498 530746 463734
rect 530982 463498 531014 463734
rect 530394 430054 531014 463498
rect 530394 429818 530426 430054
rect 530662 429818 530746 430054
rect 530982 429818 531014 430054
rect 530394 429734 531014 429818
rect 530394 429498 530426 429734
rect 530662 429498 530746 429734
rect 530982 429498 531014 429734
rect 530394 396054 531014 429498
rect 530394 395818 530426 396054
rect 530662 395818 530746 396054
rect 530982 395818 531014 396054
rect 530394 395734 531014 395818
rect 530394 395498 530426 395734
rect 530662 395498 530746 395734
rect 530982 395498 531014 395734
rect 530394 362054 531014 395498
rect 530394 361818 530426 362054
rect 530662 361818 530746 362054
rect 530982 361818 531014 362054
rect 530394 361734 531014 361818
rect 530394 361498 530426 361734
rect 530662 361498 530746 361734
rect 530982 361498 531014 361734
rect 530394 328054 531014 361498
rect 530394 327818 530426 328054
rect 530662 327818 530746 328054
rect 530982 327818 531014 328054
rect 530394 327734 531014 327818
rect 530394 327498 530426 327734
rect 530662 327498 530746 327734
rect 530982 327498 531014 327734
rect 530394 294054 531014 327498
rect 530394 293818 530426 294054
rect 530662 293818 530746 294054
rect 530982 293818 531014 294054
rect 530394 293734 531014 293818
rect 530394 293498 530426 293734
rect 530662 293498 530746 293734
rect 530982 293498 531014 293734
rect 530394 260054 531014 293498
rect 530394 259818 530426 260054
rect 530662 259818 530746 260054
rect 530982 259818 531014 260054
rect 530394 259734 531014 259818
rect 530394 259498 530426 259734
rect 530662 259498 530746 259734
rect 530982 259498 531014 259734
rect 530394 226054 531014 259498
rect 530394 225818 530426 226054
rect 530662 225818 530746 226054
rect 530982 225818 531014 226054
rect 530394 225734 531014 225818
rect 530394 225498 530426 225734
rect 530662 225498 530746 225734
rect 530982 225498 531014 225734
rect 530394 192054 531014 225498
rect 530394 191818 530426 192054
rect 530662 191818 530746 192054
rect 530982 191818 531014 192054
rect 530394 191734 531014 191818
rect 530394 191498 530426 191734
rect 530662 191498 530746 191734
rect 530982 191498 531014 191734
rect 530394 158054 531014 191498
rect 530394 157818 530426 158054
rect 530662 157818 530746 158054
rect 530982 157818 531014 158054
rect 530394 157734 531014 157818
rect 530394 157498 530426 157734
rect 530662 157498 530746 157734
rect 530982 157498 531014 157734
rect 530394 124054 531014 157498
rect 530394 123818 530426 124054
rect 530662 123818 530746 124054
rect 530982 123818 531014 124054
rect 530394 123734 531014 123818
rect 530394 123498 530426 123734
rect 530662 123498 530746 123734
rect 530982 123498 531014 123734
rect 530394 90054 531014 123498
rect 530394 89818 530426 90054
rect 530662 89818 530746 90054
rect 530982 89818 531014 90054
rect 530394 89734 531014 89818
rect 530394 89498 530426 89734
rect 530662 89498 530746 89734
rect 530982 89498 531014 89734
rect 530394 56054 531014 89498
rect 530394 55818 530426 56054
rect 530662 55818 530746 56054
rect 530982 55818 531014 56054
rect 530394 55734 531014 55818
rect 530394 55498 530426 55734
rect 530662 55498 530746 55734
rect 530982 55498 531014 55734
rect 530394 22054 531014 55498
rect 530394 21818 530426 22054
rect 530662 21818 530746 22054
rect 530982 21818 531014 22054
rect 530394 21734 531014 21818
rect 530394 21498 530426 21734
rect 530662 21498 530746 21734
rect 530982 21498 531014 21734
rect 530394 -5146 531014 21498
rect 530394 -5382 530426 -5146
rect 530662 -5382 530746 -5146
rect 530982 -5382 531014 -5146
rect 530394 -5466 531014 -5382
rect 530394 -5702 530426 -5466
rect 530662 -5702 530746 -5466
rect 530982 -5702 531014 -5466
rect 530394 -7654 531014 -5702
rect 534114 710598 534734 711590
rect 534114 710362 534146 710598
rect 534382 710362 534466 710598
rect 534702 710362 534734 710598
rect 534114 710278 534734 710362
rect 534114 710042 534146 710278
rect 534382 710042 534466 710278
rect 534702 710042 534734 710278
rect 534114 671774 534734 710042
rect 534114 671538 534146 671774
rect 534382 671538 534466 671774
rect 534702 671538 534734 671774
rect 534114 671454 534734 671538
rect 534114 671218 534146 671454
rect 534382 671218 534466 671454
rect 534702 671218 534734 671454
rect 534114 637774 534734 671218
rect 534114 637538 534146 637774
rect 534382 637538 534466 637774
rect 534702 637538 534734 637774
rect 534114 637454 534734 637538
rect 534114 637218 534146 637454
rect 534382 637218 534466 637454
rect 534702 637218 534734 637454
rect 534114 603774 534734 637218
rect 534114 603538 534146 603774
rect 534382 603538 534466 603774
rect 534702 603538 534734 603774
rect 534114 603454 534734 603538
rect 534114 603218 534146 603454
rect 534382 603218 534466 603454
rect 534702 603218 534734 603454
rect 534114 569774 534734 603218
rect 534114 569538 534146 569774
rect 534382 569538 534466 569774
rect 534702 569538 534734 569774
rect 534114 569454 534734 569538
rect 534114 569218 534146 569454
rect 534382 569218 534466 569454
rect 534702 569218 534734 569454
rect 534114 535774 534734 569218
rect 534114 535538 534146 535774
rect 534382 535538 534466 535774
rect 534702 535538 534734 535774
rect 534114 535454 534734 535538
rect 534114 535218 534146 535454
rect 534382 535218 534466 535454
rect 534702 535218 534734 535454
rect 534114 501774 534734 535218
rect 534114 501538 534146 501774
rect 534382 501538 534466 501774
rect 534702 501538 534734 501774
rect 534114 501454 534734 501538
rect 534114 501218 534146 501454
rect 534382 501218 534466 501454
rect 534702 501218 534734 501454
rect 534114 467774 534734 501218
rect 534114 467538 534146 467774
rect 534382 467538 534466 467774
rect 534702 467538 534734 467774
rect 534114 467454 534734 467538
rect 534114 467218 534146 467454
rect 534382 467218 534466 467454
rect 534702 467218 534734 467454
rect 534114 433774 534734 467218
rect 534114 433538 534146 433774
rect 534382 433538 534466 433774
rect 534702 433538 534734 433774
rect 534114 433454 534734 433538
rect 534114 433218 534146 433454
rect 534382 433218 534466 433454
rect 534702 433218 534734 433454
rect 534114 399774 534734 433218
rect 534114 399538 534146 399774
rect 534382 399538 534466 399774
rect 534702 399538 534734 399774
rect 534114 399454 534734 399538
rect 534114 399218 534146 399454
rect 534382 399218 534466 399454
rect 534702 399218 534734 399454
rect 534114 365774 534734 399218
rect 534114 365538 534146 365774
rect 534382 365538 534466 365774
rect 534702 365538 534734 365774
rect 534114 365454 534734 365538
rect 534114 365218 534146 365454
rect 534382 365218 534466 365454
rect 534702 365218 534734 365454
rect 534114 331774 534734 365218
rect 534114 331538 534146 331774
rect 534382 331538 534466 331774
rect 534702 331538 534734 331774
rect 534114 331454 534734 331538
rect 534114 331218 534146 331454
rect 534382 331218 534466 331454
rect 534702 331218 534734 331454
rect 534114 297774 534734 331218
rect 534114 297538 534146 297774
rect 534382 297538 534466 297774
rect 534702 297538 534734 297774
rect 534114 297454 534734 297538
rect 534114 297218 534146 297454
rect 534382 297218 534466 297454
rect 534702 297218 534734 297454
rect 534114 263774 534734 297218
rect 534114 263538 534146 263774
rect 534382 263538 534466 263774
rect 534702 263538 534734 263774
rect 534114 263454 534734 263538
rect 534114 263218 534146 263454
rect 534382 263218 534466 263454
rect 534702 263218 534734 263454
rect 534114 229774 534734 263218
rect 534114 229538 534146 229774
rect 534382 229538 534466 229774
rect 534702 229538 534734 229774
rect 534114 229454 534734 229538
rect 534114 229218 534146 229454
rect 534382 229218 534466 229454
rect 534702 229218 534734 229454
rect 534114 195774 534734 229218
rect 534114 195538 534146 195774
rect 534382 195538 534466 195774
rect 534702 195538 534734 195774
rect 534114 195454 534734 195538
rect 534114 195218 534146 195454
rect 534382 195218 534466 195454
rect 534702 195218 534734 195454
rect 534114 161774 534734 195218
rect 534114 161538 534146 161774
rect 534382 161538 534466 161774
rect 534702 161538 534734 161774
rect 534114 161454 534734 161538
rect 534114 161218 534146 161454
rect 534382 161218 534466 161454
rect 534702 161218 534734 161454
rect 534114 127774 534734 161218
rect 534114 127538 534146 127774
rect 534382 127538 534466 127774
rect 534702 127538 534734 127774
rect 534114 127454 534734 127538
rect 534114 127218 534146 127454
rect 534382 127218 534466 127454
rect 534702 127218 534734 127454
rect 534114 93774 534734 127218
rect 534114 93538 534146 93774
rect 534382 93538 534466 93774
rect 534702 93538 534734 93774
rect 534114 93454 534734 93538
rect 534114 93218 534146 93454
rect 534382 93218 534466 93454
rect 534702 93218 534734 93454
rect 534114 59774 534734 93218
rect 534114 59538 534146 59774
rect 534382 59538 534466 59774
rect 534702 59538 534734 59774
rect 534114 59454 534734 59538
rect 534114 59218 534146 59454
rect 534382 59218 534466 59454
rect 534702 59218 534734 59454
rect 534114 25774 534734 59218
rect 534114 25538 534146 25774
rect 534382 25538 534466 25774
rect 534702 25538 534734 25774
rect 534114 25454 534734 25538
rect 534114 25218 534146 25454
rect 534382 25218 534466 25454
rect 534702 25218 534734 25454
rect 534114 -6106 534734 25218
rect 534114 -6342 534146 -6106
rect 534382 -6342 534466 -6106
rect 534702 -6342 534734 -6106
rect 534114 -6426 534734 -6342
rect 534114 -6662 534146 -6426
rect 534382 -6662 534466 -6426
rect 534702 -6662 534734 -6426
rect 534114 -7654 534734 -6662
rect 537834 711558 538454 711590
rect 537834 711322 537866 711558
rect 538102 711322 538186 711558
rect 538422 711322 538454 711558
rect 537834 711238 538454 711322
rect 537834 711002 537866 711238
rect 538102 711002 538186 711238
rect 538422 711002 538454 711238
rect 537834 675494 538454 711002
rect 537834 675258 537866 675494
rect 538102 675258 538186 675494
rect 538422 675258 538454 675494
rect 537834 675174 538454 675258
rect 537834 674938 537866 675174
rect 538102 674938 538186 675174
rect 538422 674938 538454 675174
rect 537834 641494 538454 674938
rect 537834 641258 537866 641494
rect 538102 641258 538186 641494
rect 538422 641258 538454 641494
rect 537834 641174 538454 641258
rect 537834 640938 537866 641174
rect 538102 640938 538186 641174
rect 538422 640938 538454 641174
rect 537834 607494 538454 640938
rect 537834 607258 537866 607494
rect 538102 607258 538186 607494
rect 538422 607258 538454 607494
rect 537834 607174 538454 607258
rect 537834 606938 537866 607174
rect 538102 606938 538186 607174
rect 538422 606938 538454 607174
rect 537834 573494 538454 606938
rect 537834 573258 537866 573494
rect 538102 573258 538186 573494
rect 538422 573258 538454 573494
rect 537834 573174 538454 573258
rect 537834 572938 537866 573174
rect 538102 572938 538186 573174
rect 538422 572938 538454 573174
rect 537834 539494 538454 572938
rect 537834 539258 537866 539494
rect 538102 539258 538186 539494
rect 538422 539258 538454 539494
rect 537834 539174 538454 539258
rect 537834 538938 537866 539174
rect 538102 538938 538186 539174
rect 538422 538938 538454 539174
rect 537834 505494 538454 538938
rect 537834 505258 537866 505494
rect 538102 505258 538186 505494
rect 538422 505258 538454 505494
rect 537834 505174 538454 505258
rect 537834 504938 537866 505174
rect 538102 504938 538186 505174
rect 538422 504938 538454 505174
rect 537834 471494 538454 504938
rect 537834 471258 537866 471494
rect 538102 471258 538186 471494
rect 538422 471258 538454 471494
rect 537834 471174 538454 471258
rect 537834 470938 537866 471174
rect 538102 470938 538186 471174
rect 538422 470938 538454 471174
rect 537834 437494 538454 470938
rect 537834 437258 537866 437494
rect 538102 437258 538186 437494
rect 538422 437258 538454 437494
rect 537834 437174 538454 437258
rect 537834 436938 537866 437174
rect 538102 436938 538186 437174
rect 538422 436938 538454 437174
rect 537834 403494 538454 436938
rect 537834 403258 537866 403494
rect 538102 403258 538186 403494
rect 538422 403258 538454 403494
rect 537834 403174 538454 403258
rect 537834 402938 537866 403174
rect 538102 402938 538186 403174
rect 538422 402938 538454 403174
rect 537834 369494 538454 402938
rect 537834 369258 537866 369494
rect 538102 369258 538186 369494
rect 538422 369258 538454 369494
rect 537834 369174 538454 369258
rect 537834 368938 537866 369174
rect 538102 368938 538186 369174
rect 538422 368938 538454 369174
rect 537834 335494 538454 368938
rect 537834 335258 537866 335494
rect 538102 335258 538186 335494
rect 538422 335258 538454 335494
rect 537834 335174 538454 335258
rect 537834 334938 537866 335174
rect 538102 334938 538186 335174
rect 538422 334938 538454 335174
rect 537834 301494 538454 334938
rect 537834 301258 537866 301494
rect 538102 301258 538186 301494
rect 538422 301258 538454 301494
rect 537834 301174 538454 301258
rect 537834 300938 537866 301174
rect 538102 300938 538186 301174
rect 538422 300938 538454 301174
rect 537834 267494 538454 300938
rect 537834 267258 537866 267494
rect 538102 267258 538186 267494
rect 538422 267258 538454 267494
rect 537834 267174 538454 267258
rect 537834 266938 537866 267174
rect 538102 266938 538186 267174
rect 538422 266938 538454 267174
rect 537834 233494 538454 266938
rect 537834 233258 537866 233494
rect 538102 233258 538186 233494
rect 538422 233258 538454 233494
rect 537834 233174 538454 233258
rect 537834 232938 537866 233174
rect 538102 232938 538186 233174
rect 538422 232938 538454 233174
rect 537834 199494 538454 232938
rect 537834 199258 537866 199494
rect 538102 199258 538186 199494
rect 538422 199258 538454 199494
rect 537834 199174 538454 199258
rect 537834 198938 537866 199174
rect 538102 198938 538186 199174
rect 538422 198938 538454 199174
rect 537834 165494 538454 198938
rect 537834 165258 537866 165494
rect 538102 165258 538186 165494
rect 538422 165258 538454 165494
rect 537834 165174 538454 165258
rect 537834 164938 537866 165174
rect 538102 164938 538186 165174
rect 538422 164938 538454 165174
rect 537834 131494 538454 164938
rect 537834 131258 537866 131494
rect 538102 131258 538186 131494
rect 538422 131258 538454 131494
rect 537834 131174 538454 131258
rect 537834 130938 537866 131174
rect 538102 130938 538186 131174
rect 538422 130938 538454 131174
rect 537834 97494 538454 130938
rect 537834 97258 537866 97494
rect 538102 97258 538186 97494
rect 538422 97258 538454 97494
rect 537834 97174 538454 97258
rect 537834 96938 537866 97174
rect 538102 96938 538186 97174
rect 538422 96938 538454 97174
rect 537834 63494 538454 96938
rect 537834 63258 537866 63494
rect 538102 63258 538186 63494
rect 538422 63258 538454 63494
rect 537834 63174 538454 63258
rect 537834 62938 537866 63174
rect 538102 62938 538186 63174
rect 538422 62938 538454 63174
rect 537834 29494 538454 62938
rect 537834 29258 537866 29494
rect 538102 29258 538186 29494
rect 538422 29258 538454 29494
rect 537834 29174 538454 29258
rect 537834 28938 537866 29174
rect 538102 28938 538186 29174
rect 538422 28938 538454 29174
rect 537834 -7066 538454 28938
rect 537834 -7302 537866 -7066
rect 538102 -7302 538186 -7066
rect 538422 -7302 538454 -7066
rect 537834 -7386 538454 -7302
rect 537834 -7622 537866 -7386
rect 538102 -7622 538186 -7386
rect 538422 -7622 538454 -7386
rect 537834 -7654 538454 -7622
rect 545794 704838 546414 711590
rect 545794 704602 545826 704838
rect 546062 704602 546146 704838
rect 546382 704602 546414 704838
rect 545794 704518 546414 704602
rect 545794 704282 545826 704518
rect 546062 704282 546146 704518
rect 546382 704282 546414 704518
rect 545794 683454 546414 704282
rect 545794 683218 545826 683454
rect 546062 683218 546146 683454
rect 546382 683218 546414 683454
rect 545794 683134 546414 683218
rect 545794 682898 545826 683134
rect 546062 682898 546146 683134
rect 546382 682898 546414 683134
rect 545794 649454 546414 682898
rect 545794 649218 545826 649454
rect 546062 649218 546146 649454
rect 546382 649218 546414 649454
rect 545794 649134 546414 649218
rect 545794 648898 545826 649134
rect 546062 648898 546146 649134
rect 546382 648898 546414 649134
rect 545794 615454 546414 648898
rect 545794 615218 545826 615454
rect 546062 615218 546146 615454
rect 546382 615218 546414 615454
rect 545794 615134 546414 615218
rect 545794 614898 545826 615134
rect 546062 614898 546146 615134
rect 546382 614898 546414 615134
rect 545794 581454 546414 614898
rect 545794 581218 545826 581454
rect 546062 581218 546146 581454
rect 546382 581218 546414 581454
rect 545794 581134 546414 581218
rect 545794 580898 545826 581134
rect 546062 580898 546146 581134
rect 546382 580898 546414 581134
rect 545794 547454 546414 580898
rect 545794 547218 545826 547454
rect 546062 547218 546146 547454
rect 546382 547218 546414 547454
rect 545794 547134 546414 547218
rect 545794 546898 545826 547134
rect 546062 546898 546146 547134
rect 546382 546898 546414 547134
rect 545794 513454 546414 546898
rect 545794 513218 545826 513454
rect 546062 513218 546146 513454
rect 546382 513218 546414 513454
rect 545794 513134 546414 513218
rect 545794 512898 545826 513134
rect 546062 512898 546146 513134
rect 546382 512898 546414 513134
rect 545794 479454 546414 512898
rect 545794 479218 545826 479454
rect 546062 479218 546146 479454
rect 546382 479218 546414 479454
rect 545794 479134 546414 479218
rect 545794 478898 545826 479134
rect 546062 478898 546146 479134
rect 546382 478898 546414 479134
rect 545794 445454 546414 478898
rect 545794 445218 545826 445454
rect 546062 445218 546146 445454
rect 546382 445218 546414 445454
rect 545794 445134 546414 445218
rect 545794 444898 545826 445134
rect 546062 444898 546146 445134
rect 546382 444898 546414 445134
rect 545794 411454 546414 444898
rect 545794 411218 545826 411454
rect 546062 411218 546146 411454
rect 546382 411218 546414 411454
rect 545794 411134 546414 411218
rect 545794 410898 545826 411134
rect 546062 410898 546146 411134
rect 546382 410898 546414 411134
rect 545794 377454 546414 410898
rect 545794 377218 545826 377454
rect 546062 377218 546146 377454
rect 546382 377218 546414 377454
rect 545794 377134 546414 377218
rect 545794 376898 545826 377134
rect 546062 376898 546146 377134
rect 546382 376898 546414 377134
rect 545794 343454 546414 376898
rect 545794 343218 545826 343454
rect 546062 343218 546146 343454
rect 546382 343218 546414 343454
rect 545794 343134 546414 343218
rect 545794 342898 545826 343134
rect 546062 342898 546146 343134
rect 546382 342898 546414 343134
rect 545794 309454 546414 342898
rect 545794 309218 545826 309454
rect 546062 309218 546146 309454
rect 546382 309218 546414 309454
rect 545794 309134 546414 309218
rect 545794 308898 545826 309134
rect 546062 308898 546146 309134
rect 546382 308898 546414 309134
rect 545794 275454 546414 308898
rect 545794 275218 545826 275454
rect 546062 275218 546146 275454
rect 546382 275218 546414 275454
rect 545794 275134 546414 275218
rect 545794 274898 545826 275134
rect 546062 274898 546146 275134
rect 546382 274898 546414 275134
rect 545794 241454 546414 274898
rect 545794 241218 545826 241454
rect 546062 241218 546146 241454
rect 546382 241218 546414 241454
rect 545794 241134 546414 241218
rect 545794 240898 545826 241134
rect 546062 240898 546146 241134
rect 546382 240898 546414 241134
rect 545794 207454 546414 240898
rect 545794 207218 545826 207454
rect 546062 207218 546146 207454
rect 546382 207218 546414 207454
rect 545794 207134 546414 207218
rect 545794 206898 545826 207134
rect 546062 206898 546146 207134
rect 546382 206898 546414 207134
rect 545794 173454 546414 206898
rect 545794 173218 545826 173454
rect 546062 173218 546146 173454
rect 546382 173218 546414 173454
rect 545794 173134 546414 173218
rect 545794 172898 545826 173134
rect 546062 172898 546146 173134
rect 546382 172898 546414 173134
rect 545794 139454 546414 172898
rect 545794 139218 545826 139454
rect 546062 139218 546146 139454
rect 546382 139218 546414 139454
rect 545794 139134 546414 139218
rect 545794 138898 545826 139134
rect 546062 138898 546146 139134
rect 546382 138898 546414 139134
rect 545794 105454 546414 138898
rect 545794 105218 545826 105454
rect 546062 105218 546146 105454
rect 546382 105218 546414 105454
rect 545794 105134 546414 105218
rect 545794 104898 545826 105134
rect 546062 104898 546146 105134
rect 546382 104898 546414 105134
rect 545794 71454 546414 104898
rect 545794 71218 545826 71454
rect 546062 71218 546146 71454
rect 546382 71218 546414 71454
rect 545794 71134 546414 71218
rect 545794 70898 545826 71134
rect 546062 70898 546146 71134
rect 546382 70898 546414 71134
rect 545794 37454 546414 70898
rect 545794 37218 545826 37454
rect 546062 37218 546146 37454
rect 546382 37218 546414 37454
rect 545794 37134 546414 37218
rect 545794 36898 545826 37134
rect 546062 36898 546146 37134
rect 546382 36898 546414 37134
rect 545794 3454 546414 36898
rect 545794 3218 545826 3454
rect 546062 3218 546146 3454
rect 546382 3218 546414 3454
rect 545794 3134 546414 3218
rect 545794 2898 545826 3134
rect 546062 2898 546146 3134
rect 546382 2898 546414 3134
rect 545794 -346 546414 2898
rect 545794 -582 545826 -346
rect 546062 -582 546146 -346
rect 546382 -582 546414 -346
rect 545794 -666 546414 -582
rect 545794 -902 545826 -666
rect 546062 -902 546146 -666
rect 546382 -902 546414 -666
rect 545794 -7654 546414 -902
rect 549514 705798 550134 711590
rect 549514 705562 549546 705798
rect 549782 705562 549866 705798
rect 550102 705562 550134 705798
rect 549514 705478 550134 705562
rect 549514 705242 549546 705478
rect 549782 705242 549866 705478
rect 550102 705242 550134 705478
rect 549514 687174 550134 705242
rect 549514 686938 549546 687174
rect 549782 686938 549866 687174
rect 550102 686938 550134 687174
rect 549514 686854 550134 686938
rect 549514 686618 549546 686854
rect 549782 686618 549866 686854
rect 550102 686618 550134 686854
rect 549514 653174 550134 686618
rect 549514 652938 549546 653174
rect 549782 652938 549866 653174
rect 550102 652938 550134 653174
rect 549514 652854 550134 652938
rect 549514 652618 549546 652854
rect 549782 652618 549866 652854
rect 550102 652618 550134 652854
rect 549514 619174 550134 652618
rect 549514 618938 549546 619174
rect 549782 618938 549866 619174
rect 550102 618938 550134 619174
rect 549514 618854 550134 618938
rect 549514 618618 549546 618854
rect 549782 618618 549866 618854
rect 550102 618618 550134 618854
rect 549514 585174 550134 618618
rect 549514 584938 549546 585174
rect 549782 584938 549866 585174
rect 550102 584938 550134 585174
rect 549514 584854 550134 584938
rect 549514 584618 549546 584854
rect 549782 584618 549866 584854
rect 550102 584618 550134 584854
rect 549514 551174 550134 584618
rect 549514 550938 549546 551174
rect 549782 550938 549866 551174
rect 550102 550938 550134 551174
rect 549514 550854 550134 550938
rect 549514 550618 549546 550854
rect 549782 550618 549866 550854
rect 550102 550618 550134 550854
rect 549514 517174 550134 550618
rect 549514 516938 549546 517174
rect 549782 516938 549866 517174
rect 550102 516938 550134 517174
rect 549514 516854 550134 516938
rect 549514 516618 549546 516854
rect 549782 516618 549866 516854
rect 550102 516618 550134 516854
rect 549514 483174 550134 516618
rect 549514 482938 549546 483174
rect 549782 482938 549866 483174
rect 550102 482938 550134 483174
rect 549514 482854 550134 482938
rect 549514 482618 549546 482854
rect 549782 482618 549866 482854
rect 550102 482618 550134 482854
rect 549514 449174 550134 482618
rect 549514 448938 549546 449174
rect 549782 448938 549866 449174
rect 550102 448938 550134 449174
rect 549514 448854 550134 448938
rect 549514 448618 549546 448854
rect 549782 448618 549866 448854
rect 550102 448618 550134 448854
rect 549514 415174 550134 448618
rect 549514 414938 549546 415174
rect 549782 414938 549866 415174
rect 550102 414938 550134 415174
rect 549514 414854 550134 414938
rect 549514 414618 549546 414854
rect 549782 414618 549866 414854
rect 550102 414618 550134 414854
rect 549514 381174 550134 414618
rect 549514 380938 549546 381174
rect 549782 380938 549866 381174
rect 550102 380938 550134 381174
rect 549514 380854 550134 380938
rect 549514 380618 549546 380854
rect 549782 380618 549866 380854
rect 550102 380618 550134 380854
rect 549514 347174 550134 380618
rect 549514 346938 549546 347174
rect 549782 346938 549866 347174
rect 550102 346938 550134 347174
rect 549514 346854 550134 346938
rect 549514 346618 549546 346854
rect 549782 346618 549866 346854
rect 550102 346618 550134 346854
rect 549514 313174 550134 346618
rect 549514 312938 549546 313174
rect 549782 312938 549866 313174
rect 550102 312938 550134 313174
rect 549514 312854 550134 312938
rect 549514 312618 549546 312854
rect 549782 312618 549866 312854
rect 550102 312618 550134 312854
rect 549514 279174 550134 312618
rect 549514 278938 549546 279174
rect 549782 278938 549866 279174
rect 550102 278938 550134 279174
rect 549514 278854 550134 278938
rect 549514 278618 549546 278854
rect 549782 278618 549866 278854
rect 550102 278618 550134 278854
rect 549514 245174 550134 278618
rect 549514 244938 549546 245174
rect 549782 244938 549866 245174
rect 550102 244938 550134 245174
rect 549514 244854 550134 244938
rect 549514 244618 549546 244854
rect 549782 244618 549866 244854
rect 550102 244618 550134 244854
rect 549514 211174 550134 244618
rect 549514 210938 549546 211174
rect 549782 210938 549866 211174
rect 550102 210938 550134 211174
rect 549514 210854 550134 210938
rect 549514 210618 549546 210854
rect 549782 210618 549866 210854
rect 550102 210618 550134 210854
rect 549514 177174 550134 210618
rect 549514 176938 549546 177174
rect 549782 176938 549866 177174
rect 550102 176938 550134 177174
rect 549514 176854 550134 176938
rect 549514 176618 549546 176854
rect 549782 176618 549866 176854
rect 550102 176618 550134 176854
rect 549514 143174 550134 176618
rect 549514 142938 549546 143174
rect 549782 142938 549866 143174
rect 550102 142938 550134 143174
rect 549514 142854 550134 142938
rect 549514 142618 549546 142854
rect 549782 142618 549866 142854
rect 550102 142618 550134 142854
rect 549514 109174 550134 142618
rect 549514 108938 549546 109174
rect 549782 108938 549866 109174
rect 550102 108938 550134 109174
rect 549514 108854 550134 108938
rect 549514 108618 549546 108854
rect 549782 108618 549866 108854
rect 550102 108618 550134 108854
rect 549514 75174 550134 108618
rect 549514 74938 549546 75174
rect 549782 74938 549866 75174
rect 550102 74938 550134 75174
rect 549514 74854 550134 74938
rect 549514 74618 549546 74854
rect 549782 74618 549866 74854
rect 550102 74618 550134 74854
rect 549514 41174 550134 74618
rect 549514 40938 549546 41174
rect 549782 40938 549866 41174
rect 550102 40938 550134 41174
rect 549514 40854 550134 40938
rect 549514 40618 549546 40854
rect 549782 40618 549866 40854
rect 550102 40618 550134 40854
rect 549514 7174 550134 40618
rect 549514 6938 549546 7174
rect 549782 6938 549866 7174
rect 550102 6938 550134 7174
rect 549514 6854 550134 6938
rect 549514 6618 549546 6854
rect 549782 6618 549866 6854
rect 550102 6618 550134 6854
rect 549514 -1306 550134 6618
rect 549514 -1542 549546 -1306
rect 549782 -1542 549866 -1306
rect 550102 -1542 550134 -1306
rect 549514 -1626 550134 -1542
rect 549514 -1862 549546 -1626
rect 549782 -1862 549866 -1626
rect 550102 -1862 550134 -1626
rect 549514 -7654 550134 -1862
rect 553234 706758 553854 711590
rect 553234 706522 553266 706758
rect 553502 706522 553586 706758
rect 553822 706522 553854 706758
rect 553234 706438 553854 706522
rect 553234 706202 553266 706438
rect 553502 706202 553586 706438
rect 553822 706202 553854 706438
rect 553234 690894 553854 706202
rect 553234 690658 553266 690894
rect 553502 690658 553586 690894
rect 553822 690658 553854 690894
rect 553234 690574 553854 690658
rect 553234 690338 553266 690574
rect 553502 690338 553586 690574
rect 553822 690338 553854 690574
rect 553234 656894 553854 690338
rect 553234 656658 553266 656894
rect 553502 656658 553586 656894
rect 553822 656658 553854 656894
rect 553234 656574 553854 656658
rect 553234 656338 553266 656574
rect 553502 656338 553586 656574
rect 553822 656338 553854 656574
rect 553234 622894 553854 656338
rect 553234 622658 553266 622894
rect 553502 622658 553586 622894
rect 553822 622658 553854 622894
rect 553234 622574 553854 622658
rect 553234 622338 553266 622574
rect 553502 622338 553586 622574
rect 553822 622338 553854 622574
rect 553234 588894 553854 622338
rect 553234 588658 553266 588894
rect 553502 588658 553586 588894
rect 553822 588658 553854 588894
rect 553234 588574 553854 588658
rect 553234 588338 553266 588574
rect 553502 588338 553586 588574
rect 553822 588338 553854 588574
rect 553234 554894 553854 588338
rect 553234 554658 553266 554894
rect 553502 554658 553586 554894
rect 553822 554658 553854 554894
rect 553234 554574 553854 554658
rect 553234 554338 553266 554574
rect 553502 554338 553586 554574
rect 553822 554338 553854 554574
rect 553234 520894 553854 554338
rect 553234 520658 553266 520894
rect 553502 520658 553586 520894
rect 553822 520658 553854 520894
rect 553234 520574 553854 520658
rect 553234 520338 553266 520574
rect 553502 520338 553586 520574
rect 553822 520338 553854 520574
rect 553234 486894 553854 520338
rect 553234 486658 553266 486894
rect 553502 486658 553586 486894
rect 553822 486658 553854 486894
rect 553234 486574 553854 486658
rect 553234 486338 553266 486574
rect 553502 486338 553586 486574
rect 553822 486338 553854 486574
rect 553234 452894 553854 486338
rect 553234 452658 553266 452894
rect 553502 452658 553586 452894
rect 553822 452658 553854 452894
rect 553234 452574 553854 452658
rect 553234 452338 553266 452574
rect 553502 452338 553586 452574
rect 553822 452338 553854 452574
rect 553234 418894 553854 452338
rect 553234 418658 553266 418894
rect 553502 418658 553586 418894
rect 553822 418658 553854 418894
rect 553234 418574 553854 418658
rect 553234 418338 553266 418574
rect 553502 418338 553586 418574
rect 553822 418338 553854 418574
rect 553234 384894 553854 418338
rect 553234 384658 553266 384894
rect 553502 384658 553586 384894
rect 553822 384658 553854 384894
rect 553234 384574 553854 384658
rect 553234 384338 553266 384574
rect 553502 384338 553586 384574
rect 553822 384338 553854 384574
rect 553234 350894 553854 384338
rect 553234 350658 553266 350894
rect 553502 350658 553586 350894
rect 553822 350658 553854 350894
rect 553234 350574 553854 350658
rect 553234 350338 553266 350574
rect 553502 350338 553586 350574
rect 553822 350338 553854 350574
rect 553234 316894 553854 350338
rect 553234 316658 553266 316894
rect 553502 316658 553586 316894
rect 553822 316658 553854 316894
rect 553234 316574 553854 316658
rect 553234 316338 553266 316574
rect 553502 316338 553586 316574
rect 553822 316338 553854 316574
rect 553234 282894 553854 316338
rect 553234 282658 553266 282894
rect 553502 282658 553586 282894
rect 553822 282658 553854 282894
rect 553234 282574 553854 282658
rect 553234 282338 553266 282574
rect 553502 282338 553586 282574
rect 553822 282338 553854 282574
rect 553234 248894 553854 282338
rect 553234 248658 553266 248894
rect 553502 248658 553586 248894
rect 553822 248658 553854 248894
rect 553234 248574 553854 248658
rect 553234 248338 553266 248574
rect 553502 248338 553586 248574
rect 553822 248338 553854 248574
rect 553234 214894 553854 248338
rect 553234 214658 553266 214894
rect 553502 214658 553586 214894
rect 553822 214658 553854 214894
rect 553234 214574 553854 214658
rect 553234 214338 553266 214574
rect 553502 214338 553586 214574
rect 553822 214338 553854 214574
rect 553234 180894 553854 214338
rect 553234 180658 553266 180894
rect 553502 180658 553586 180894
rect 553822 180658 553854 180894
rect 553234 180574 553854 180658
rect 553234 180338 553266 180574
rect 553502 180338 553586 180574
rect 553822 180338 553854 180574
rect 553234 146894 553854 180338
rect 553234 146658 553266 146894
rect 553502 146658 553586 146894
rect 553822 146658 553854 146894
rect 553234 146574 553854 146658
rect 553234 146338 553266 146574
rect 553502 146338 553586 146574
rect 553822 146338 553854 146574
rect 553234 112894 553854 146338
rect 553234 112658 553266 112894
rect 553502 112658 553586 112894
rect 553822 112658 553854 112894
rect 553234 112574 553854 112658
rect 553234 112338 553266 112574
rect 553502 112338 553586 112574
rect 553822 112338 553854 112574
rect 553234 78894 553854 112338
rect 553234 78658 553266 78894
rect 553502 78658 553586 78894
rect 553822 78658 553854 78894
rect 553234 78574 553854 78658
rect 553234 78338 553266 78574
rect 553502 78338 553586 78574
rect 553822 78338 553854 78574
rect 553234 44894 553854 78338
rect 553234 44658 553266 44894
rect 553502 44658 553586 44894
rect 553822 44658 553854 44894
rect 553234 44574 553854 44658
rect 553234 44338 553266 44574
rect 553502 44338 553586 44574
rect 553822 44338 553854 44574
rect 553234 10894 553854 44338
rect 553234 10658 553266 10894
rect 553502 10658 553586 10894
rect 553822 10658 553854 10894
rect 553234 10574 553854 10658
rect 553234 10338 553266 10574
rect 553502 10338 553586 10574
rect 553822 10338 553854 10574
rect 553234 -2266 553854 10338
rect 553234 -2502 553266 -2266
rect 553502 -2502 553586 -2266
rect 553822 -2502 553854 -2266
rect 553234 -2586 553854 -2502
rect 553234 -2822 553266 -2586
rect 553502 -2822 553586 -2586
rect 553822 -2822 553854 -2586
rect 553234 -7654 553854 -2822
rect 556954 707718 557574 711590
rect 556954 707482 556986 707718
rect 557222 707482 557306 707718
rect 557542 707482 557574 707718
rect 556954 707398 557574 707482
rect 556954 707162 556986 707398
rect 557222 707162 557306 707398
rect 557542 707162 557574 707398
rect 556954 694614 557574 707162
rect 556954 694378 556986 694614
rect 557222 694378 557306 694614
rect 557542 694378 557574 694614
rect 556954 694294 557574 694378
rect 556954 694058 556986 694294
rect 557222 694058 557306 694294
rect 557542 694058 557574 694294
rect 556954 660614 557574 694058
rect 556954 660378 556986 660614
rect 557222 660378 557306 660614
rect 557542 660378 557574 660614
rect 556954 660294 557574 660378
rect 556954 660058 556986 660294
rect 557222 660058 557306 660294
rect 557542 660058 557574 660294
rect 556954 626614 557574 660058
rect 556954 626378 556986 626614
rect 557222 626378 557306 626614
rect 557542 626378 557574 626614
rect 556954 626294 557574 626378
rect 556954 626058 556986 626294
rect 557222 626058 557306 626294
rect 557542 626058 557574 626294
rect 556954 592614 557574 626058
rect 556954 592378 556986 592614
rect 557222 592378 557306 592614
rect 557542 592378 557574 592614
rect 556954 592294 557574 592378
rect 556954 592058 556986 592294
rect 557222 592058 557306 592294
rect 557542 592058 557574 592294
rect 556954 558614 557574 592058
rect 556954 558378 556986 558614
rect 557222 558378 557306 558614
rect 557542 558378 557574 558614
rect 556954 558294 557574 558378
rect 556954 558058 556986 558294
rect 557222 558058 557306 558294
rect 557542 558058 557574 558294
rect 556954 524614 557574 558058
rect 556954 524378 556986 524614
rect 557222 524378 557306 524614
rect 557542 524378 557574 524614
rect 556954 524294 557574 524378
rect 556954 524058 556986 524294
rect 557222 524058 557306 524294
rect 557542 524058 557574 524294
rect 556954 490614 557574 524058
rect 556954 490378 556986 490614
rect 557222 490378 557306 490614
rect 557542 490378 557574 490614
rect 556954 490294 557574 490378
rect 556954 490058 556986 490294
rect 557222 490058 557306 490294
rect 557542 490058 557574 490294
rect 556954 456614 557574 490058
rect 556954 456378 556986 456614
rect 557222 456378 557306 456614
rect 557542 456378 557574 456614
rect 556954 456294 557574 456378
rect 556954 456058 556986 456294
rect 557222 456058 557306 456294
rect 557542 456058 557574 456294
rect 556954 422614 557574 456058
rect 556954 422378 556986 422614
rect 557222 422378 557306 422614
rect 557542 422378 557574 422614
rect 556954 422294 557574 422378
rect 556954 422058 556986 422294
rect 557222 422058 557306 422294
rect 557542 422058 557574 422294
rect 556954 388614 557574 422058
rect 556954 388378 556986 388614
rect 557222 388378 557306 388614
rect 557542 388378 557574 388614
rect 556954 388294 557574 388378
rect 556954 388058 556986 388294
rect 557222 388058 557306 388294
rect 557542 388058 557574 388294
rect 556954 354614 557574 388058
rect 556954 354378 556986 354614
rect 557222 354378 557306 354614
rect 557542 354378 557574 354614
rect 556954 354294 557574 354378
rect 556954 354058 556986 354294
rect 557222 354058 557306 354294
rect 557542 354058 557574 354294
rect 556954 320614 557574 354058
rect 556954 320378 556986 320614
rect 557222 320378 557306 320614
rect 557542 320378 557574 320614
rect 556954 320294 557574 320378
rect 556954 320058 556986 320294
rect 557222 320058 557306 320294
rect 557542 320058 557574 320294
rect 556954 286614 557574 320058
rect 556954 286378 556986 286614
rect 557222 286378 557306 286614
rect 557542 286378 557574 286614
rect 556954 286294 557574 286378
rect 556954 286058 556986 286294
rect 557222 286058 557306 286294
rect 557542 286058 557574 286294
rect 556954 252614 557574 286058
rect 556954 252378 556986 252614
rect 557222 252378 557306 252614
rect 557542 252378 557574 252614
rect 556954 252294 557574 252378
rect 556954 252058 556986 252294
rect 557222 252058 557306 252294
rect 557542 252058 557574 252294
rect 556954 218614 557574 252058
rect 556954 218378 556986 218614
rect 557222 218378 557306 218614
rect 557542 218378 557574 218614
rect 556954 218294 557574 218378
rect 556954 218058 556986 218294
rect 557222 218058 557306 218294
rect 557542 218058 557574 218294
rect 556954 184614 557574 218058
rect 556954 184378 556986 184614
rect 557222 184378 557306 184614
rect 557542 184378 557574 184614
rect 556954 184294 557574 184378
rect 556954 184058 556986 184294
rect 557222 184058 557306 184294
rect 557542 184058 557574 184294
rect 556954 150614 557574 184058
rect 556954 150378 556986 150614
rect 557222 150378 557306 150614
rect 557542 150378 557574 150614
rect 556954 150294 557574 150378
rect 556954 150058 556986 150294
rect 557222 150058 557306 150294
rect 557542 150058 557574 150294
rect 556954 116614 557574 150058
rect 556954 116378 556986 116614
rect 557222 116378 557306 116614
rect 557542 116378 557574 116614
rect 556954 116294 557574 116378
rect 556954 116058 556986 116294
rect 557222 116058 557306 116294
rect 557542 116058 557574 116294
rect 556954 82614 557574 116058
rect 556954 82378 556986 82614
rect 557222 82378 557306 82614
rect 557542 82378 557574 82614
rect 556954 82294 557574 82378
rect 556954 82058 556986 82294
rect 557222 82058 557306 82294
rect 557542 82058 557574 82294
rect 556954 48614 557574 82058
rect 556954 48378 556986 48614
rect 557222 48378 557306 48614
rect 557542 48378 557574 48614
rect 556954 48294 557574 48378
rect 556954 48058 556986 48294
rect 557222 48058 557306 48294
rect 557542 48058 557574 48294
rect 556954 14614 557574 48058
rect 556954 14378 556986 14614
rect 557222 14378 557306 14614
rect 557542 14378 557574 14614
rect 556954 14294 557574 14378
rect 556954 14058 556986 14294
rect 557222 14058 557306 14294
rect 557542 14058 557574 14294
rect 556954 -3226 557574 14058
rect 556954 -3462 556986 -3226
rect 557222 -3462 557306 -3226
rect 557542 -3462 557574 -3226
rect 556954 -3546 557574 -3462
rect 556954 -3782 556986 -3546
rect 557222 -3782 557306 -3546
rect 557542 -3782 557574 -3546
rect 556954 -7654 557574 -3782
rect 560674 708678 561294 711590
rect 560674 708442 560706 708678
rect 560942 708442 561026 708678
rect 561262 708442 561294 708678
rect 560674 708358 561294 708442
rect 560674 708122 560706 708358
rect 560942 708122 561026 708358
rect 561262 708122 561294 708358
rect 560674 698334 561294 708122
rect 560674 698098 560706 698334
rect 560942 698098 561026 698334
rect 561262 698098 561294 698334
rect 560674 698014 561294 698098
rect 560674 697778 560706 698014
rect 560942 697778 561026 698014
rect 561262 697778 561294 698014
rect 560674 664334 561294 697778
rect 560674 664098 560706 664334
rect 560942 664098 561026 664334
rect 561262 664098 561294 664334
rect 560674 664014 561294 664098
rect 560674 663778 560706 664014
rect 560942 663778 561026 664014
rect 561262 663778 561294 664014
rect 560674 630334 561294 663778
rect 560674 630098 560706 630334
rect 560942 630098 561026 630334
rect 561262 630098 561294 630334
rect 560674 630014 561294 630098
rect 560674 629778 560706 630014
rect 560942 629778 561026 630014
rect 561262 629778 561294 630014
rect 560674 596334 561294 629778
rect 560674 596098 560706 596334
rect 560942 596098 561026 596334
rect 561262 596098 561294 596334
rect 560674 596014 561294 596098
rect 560674 595778 560706 596014
rect 560942 595778 561026 596014
rect 561262 595778 561294 596014
rect 560674 562334 561294 595778
rect 560674 562098 560706 562334
rect 560942 562098 561026 562334
rect 561262 562098 561294 562334
rect 560674 562014 561294 562098
rect 560674 561778 560706 562014
rect 560942 561778 561026 562014
rect 561262 561778 561294 562014
rect 560674 528334 561294 561778
rect 560674 528098 560706 528334
rect 560942 528098 561026 528334
rect 561262 528098 561294 528334
rect 560674 528014 561294 528098
rect 560674 527778 560706 528014
rect 560942 527778 561026 528014
rect 561262 527778 561294 528014
rect 560674 494334 561294 527778
rect 560674 494098 560706 494334
rect 560942 494098 561026 494334
rect 561262 494098 561294 494334
rect 560674 494014 561294 494098
rect 560674 493778 560706 494014
rect 560942 493778 561026 494014
rect 561262 493778 561294 494014
rect 560674 460334 561294 493778
rect 560674 460098 560706 460334
rect 560942 460098 561026 460334
rect 561262 460098 561294 460334
rect 560674 460014 561294 460098
rect 560674 459778 560706 460014
rect 560942 459778 561026 460014
rect 561262 459778 561294 460014
rect 560674 426334 561294 459778
rect 560674 426098 560706 426334
rect 560942 426098 561026 426334
rect 561262 426098 561294 426334
rect 560674 426014 561294 426098
rect 560674 425778 560706 426014
rect 560942 425778 561026 426014
rect 561262 425778 561294 426014
rect 560674 392334 561294 425778
rect 560674 392098 560706 392334
rect 560942 392098 561026 392334
rect 561262 392098 561294 392334
rect 560674 392014 561294 392098
rect 560674 391778 560706 392014
rect 560942 391778 561026 392014
rect 561262 391778 561294 392014
rect 560674 358334 561294 391778
rect 560674 358098 560706 358334
rect 560942 358098 561026 358334
rect 561262 358098 561294 358334
rect 560674 358014 561294 358098
rect 560674 357778 560706 358014
rect 560942 357778 561026 358014
rect 561262 357778 561294 358014
rect 560674 324334 561294 357778
rect 560674 324098 560706 324334
rect 560942 324098 561026 324334
rect 561262 324098 561294 324334
rect 560674 324014 561294 324098
rect 560674 323778 560706 324014
rect 560942 323778 561026 324014
rect 561262 323778 561294 324014
rect 560674 290334 561294 323778
rect 560674 290098 560706 290334
rect 560942 290098 561026 290334
rect 561262 290098 561294 290334
rect 560674 290014 561294 290098
rect 560674 289778 560706 290014
rect 560942 289778 561026 290014
rect 561262 289778 561294 290014
rect 560674 256334 561294 289778
rect 560674 256098 560706 256334
rect 560942 256098 561026 256334
rect 561262 256098 561294 256334
rect 560674 256014 561294 256098
rect 560674 255778 560706 256014
rect 560942 255778 561026 256014
rect 561262 255778 561294 256014
rect 560674 222334 561294 255778
rect 560674 222098 560706 222334
rect 560942 222098 561026 222334
rect 561262 222098 561294 222334
rect 560674 222014 561294 222098
rect 560674 221778 560706 222014
rect 560942 221778 561026 222014
rect 561262 221778 561294 222014
rect 560674 188334 561294 221778
rect 560674 188098 560706 188334
rect 560942 188098 561026 188334
rect 561262 188098 561294 188334
rect 560674 188014 561294 188098
rect 560674 187778 560706 188014
rect 560942 187778 561026 188014
rect 561262 187778 561294 188014
rect 560674 154334 561294 187778
rect 560674 154098 560706 154334
rect 560942 154098 561026 154334
rect 561262 154098 561294 154334
rect 560674 154014 561294 154098
rect 560674 153778 560706 154014
rect 560942 153778 561026 154014
rect 561262 153778 561294 154014
rect 560674 120334 561294 153778
rect 560674 120098 560706 120334
rect 560942 120098 561026 120334
rect 561262 120098 561294 120334
rect 560674 120014 561294 120098
rect 560674 119778 560706 120014
rect 560942 119778 561026 120014
rect 561262 119778 561294 120014
rect 560674 86334 561294 119778
rect 560674 86098 560706 86334
rect 560942 86098 561026 86334
rect 561262 86098 561294 86334
rect 560674 86014 561294 86098
rect 560674 85778 560706 86014
rect 560942 85778 561026 86014
rect 561262 85778 561294 86014
rect 560674 52334 561294 85778
rect 560674 52098 560706 52334
rect 560942 52098 561026 52334
rect 561262 52098 561294 52334
rect 560674 52014 561294 52098
rect 560674 51778 560706 52014
rect 560942 51778 561026 52014
rect 561262 51778 561294 52014
rect 560674 18334 561294 51778
rect 560674 18098 560706 18334
rect 560942 18098 561026 18334
rect 561262 18098 561294 18334
rect 560674 18014 561294 18098
rect 560674 17778 560706 18014
rect 560942 17778 561026 18014
rect 561262 17778 561294 18014
rect 560674 -4186 561294 17778
rect 560674 -4422 560706 -4186
rect 560942 -4422 561026 -4186
rect 561262 -4422 561294 -4186
rect 560674 -4506 561294 -4422
rect 560674 -4742 560706 -4506
rect 560942 -4742 561026 -4506
rect 561262 -4742 561294 -4506
rect 560674 -7654 561294 -4742
rect 564394 709638 565014 711590
rect 564394 709402 564426 709638
rect 564662 709402 564746 709638
rect 564982 709402 565014 709638
rect 564394 709318 565014 709402
rect 564394 709082 564426 709318
rect 564662 709082 564746 709318
rect 564982 709082 565014 709318
rect 564394 668054 565014 709082
rect 564394 667818 564426 668054
rect 564662 667818 564746 668054
rect 564982 667818 565014 668054
rect 564394 667734 565014 667818
rect 564394 667498 564426 667734
rect 564662 667498 564746 667734
rect 564982 667498 565014 667734
rect 564394 634054 565014 667498
rect 564394 633818 564426 634054
rect 564662 633818 564746 634054
rect 564982 633818 565014 634054
rect 564394 633734 565014 633818
rect 564394 633498 564426 633734
rect 564662 633498 564746 633734
rect 564982 633498 565014 633734
rect 564394 600054 565014 633498
rect 564394 599818 564426 600054
rect 564662 599818 564746 600054
rect 564982 599818 565014 600054
rect 564394 599734 565014 599818
rect 564394 599498 564426 599734
rect 564662 599498 564746 599734
rect 564982 599498 565014 599734
rect 564394 566054 565014 599498
rect 564394 565818 564426 566054
rect 564662 565818 564746 566054
rect 564982 565818 565014 566054
rect 564394 565734 565014 565818
rect 564394 565498 564426 565734
rect 564662 565498 564746 565734
rect 564982 565498 565014 565734
rect 564394 532054 565014 565498
rect 564394 531818 564426 532054
rect 564662 531818 564746 532054
rect 564982 531818 565014 532054
rect 564394 531734 565014 531818
rect 564394 531498 564426 531734
rect 564662 531498 564746 531734
rect 564982 531498 565014 531734
rect 564394 498054 565014 531498
rect 564394 497818 564426 498054
rect 564662 497818 564746 498054
rect 564982 497818 565014 498054
rect 564394 497734 565014 497818
rect 564394 497498 564426 497734
rect 564662 497498 564746 497734
rect 564982 497498 565014 497734
rect 564394 464054 565014 497498
rect 564394 463818 564426 464054
rect 564662 463818 564746 464054
rect 564982 463818 565014 464054
rect 564394 463734 565014 463818
rect 564394 463498 564426 463734
rect 564662 463498 564746 463734
rect 564982 463498 565014 463734
rect 564394 430054 565014 463498
rect 564394 429818 564426 430054
rect 564662 429818 564746 430054
rect 564982 429818 565014 430054
rect 564394 429734 565014 429818
rect 564394 429498 564426 429734
rect 564662 429498 564746 429734
rect 564982 429498 565014 429734
rect 564394 396054 565014 429498
rect 564394 395818 564426 396054
rect 564662 395818 564746 396054
rect 564982 395818 565014 396054
rect 564394 395734 565014 395818
rect 564394 395498 564426 395734
rect 564662 395498 564746 395734
rect 564982 395498 565014 395734
rect 564394 362054 565014 395498
rect 564394 361818 564426 362054
rect 564662 361818 564746 362054
rect 564982 361818 565014 362054
rect 564394 361734 565014 361818
rect 564394 361498 564426 361734
rect 564662 361498 564746 361734
rect 564982 361498 565014 361734
rect 564394 328054 565014 361498
rect 564394 327818 564426 328054
rect 564662 327818 564746 328054
rect 564982 327818 565014 328054
rect 564394 327734 565014 327818
rect 564394 327498 564426 327734
rect 564662 327498 564746 327734
rect 564982 327498 565014 327734
rect 564394 294054 565014 327498
rect 564394 293818 564426 294054
rect 564662 293818 564746 294054
rect 564982 293818 565014 294054
rect 564394 293734 565014 293818
rect 564394 293498 564426 293734
rect 564662 293498 564746 293734
rect 564982 293498 565014 293734
rect 564394 260054 565014 293498
rect 564394 259818 564426 260054
rect 564662 259818 564746 260054
rect 564982 259818 565014 260054
rect 564394 259734 565014 259818
rect 564394 259498 564426 259734
rect 564662 259498 564746 259734
rect 564982 259498 565014 259734
rect 564394 226054 565014 259498
rect 564394 225818 564426 226054
rect 564662 225818 564746 226054
rect 564982 225818 565014 226054
rect 564394 225734 565014 225818
rect 564394 225498 564426 225734
rect 564662 225498 564746 225734
rect 564982 225498 565014 225734
rect 564394 192054 565014 225498
rect 564394 191818 564426 192054
rect 564662 191818 564746 192054
rect 564982 191818 565014 192054
rect 564394 191734 565014 191818
rect 564394 191498 564426 191734
rect 564662 191498 564746 191734
rect 564982 191498 565014 191734
rect 564394 158054 565014 191498
rect 564394 157818 564426 158054
rect 564662 157818 564746 158054
rect 564982 157818 565014 158054
rect 564394 157734 565014 157818
rect 564394 157498 564426 157734
rect 564662 157498 564746 157734
rect 564982 157498 565014 157734
rect 564394 124054 565014 157498
rect 564394 123818 564426 124054
rect 564662 123818 564746 124054
rect 564982 123818 565014 124054
rect 564394 123734 565014 123818
rect 564394 123498 564426 123734
rect 564662 123498 564746 123734
rect 564982 123498 565014 123734
rect 564394 90054 565014 123498
rect 564394 89818 564426 90054
rect 564662 89818 564746 90054
rect 564982 89818 565014 90054
rect 564394 89734 565014 89818
rect 564394 89498 564426 89734
rect 564662 89498 564746 89734
rect 564982 89498 565014 89734
rect 564394 56054 565014 89498
rect 564394 55818 564426 56054
rect 564662 55818 564746 56054
rect 564982 55818 565014 56054
rect 564394 55734 565014 55818
rect 564394 55498 564426 55734
rect 564662 55498 564746 55734
rect 564982 55498 565014 55734
rect 564394 22054 565014 55498
rect 564394 21818 564426 22054
rect 564662 21818 564746 22054
rect 564982 21818 565014 22054
rect 564394 21734 565014 21818
rect 564394 21498 564426 21734
rect 564662 21498 564746 21734
rect 564982 21498 565014 21734
rect 564394 -5146 565014 21498
rect 564394 -5382 564426 -5146
rect 564662 -5382 564746 -5146
rect 564982 -5382 565014 -5146
rect 564394 -5466 565014 -5382
rect 564394 -5702 564426 -5466
rect 564662 -5702 564746 -5466
rect 564982 -5702 565014 -5466
rect 564394 -7654 565014 -5702
rect 568114 710598 568734 711590
rect 568114 710362 568146 710598
rect 568382 710362 568466 710598
rect 568702 710362 568734 710598
rect 568114 710278 568734 710362
rect 568114 710042 568146 710278
rect 568382 710042 568466 710278
rect 568702 710042 568734 710278
rect 568114 671774 568734 710042
rect 568114 671538 568146 671774
rect 568382 671538 568466 671774
rect 568702 671538 568734 671774
rect 568114 671454 568734 671538
rect 568114 671218 568146 671454
rect 568382 671218 568466 671454
rect 568702 671218 568734 671454
rect 568114 637774 568734 671218
rect 568114 637538 568146 637774
rect 568382 637538 568466 637774
rect 568702 637538 568734 637774
rect 568114 637454 568734 637538
rect 568114 637218 568146 637454
rect 568382 637218 568466 637454
rect 568702 637218 568734 637454
rect 568114 603774 568734 637218
rect 568114 603538 568146 603774
rect 568382 603538 568466 603774
rect 568702 603538 568734 603774
rect 568114 603454 568734 603538
rect 568114 603218 568146 603454
rect 568382 603218 568466 603454
rect 568702 603218 568734 603454
rect 568114 569774 568734 603218
rect 568114 569538 568146 569774
rect 568382 569538 568466 569774
rect 568702 569538 568734 569774
rect 568114 569454 568734 569538
rect 568114 569218 568146 569454
rect 568382 569218 568466 569454
rect 568702 569218 568734 569454
rect 568114 535774 568734 569218
rect 568114 535538 568146 535774
rect 568382 535538 568466 535774
rect 568702 535538 568734 535774
rect 568114 535454 568734 535538
rect 568114 535218 568146 535454
rect 568382 535218 568466 535454
rect 568702 535218 568734 535454
rect 568114 501774 568734 535218
rect 568114 501538 568146 501774
rect 568382 501538 568466 501774
rect 568702 501538 568734 501774
rect 568114 501454 568734 501538
rect 568114 501218 568146 501454
rect 568382 501218 568466 501454
rect 568702 501218 568734 501454
rect 568114 467774 568734 501218
rect 568114 467538 568146 467774
rect 568382 467538 568466 467774
rect 568702 467538 568734 467774
rect 568114 467454 568734 467538
rect 568114 467218 568146 467454
rect 568382 467218 568466 467454
rect 568702 467218 568734 467454
rect 568114 433774 568734 467218
rect 568114 433538 568146 433774
rect 568382 433538 568466 433774
rect 568702 433538 568734 433774
rect 568114 433454 568734 433538
rect 568114 433218 568146 433454
rect 568382 433218 568466 433454
rect 568702 433218 568734 433454
rect 568114 399774 568734 433218
rect 568114 399538 568146 399774
rect 568382 399538 568466 399774
rect 568702 399538 568734 399774
rect 568114 399454 568734 399538
rect 568114 399218 568146 399454
rect 568382 399218 568466 399454
rect 568702 399218 568734 399454
rect 568114 365774 568734 399218
rect 568114 365538 568146 365774
rect 568382 365538 568466 365774
rect 568702 365538 568734 365774
rect 568114 365454 568734 365538
rect 568114 365218 568146 365454
rect 568382 365218 568466 365454
rect 568702 365218 568734 365454
rect 568114 331774 568734 365218
rect 568114 331538 568146 331774
rect 568382 331538 568466 331774
rect 568702 331538 568734 331774
rect 568114 331454 568734 331538
rect 568114 331218 568146 331454
rect 568382 331218 568466 331454
rect 568702 331218 568734 331454
rect 568114 297774 568734 331218
rect 568114 297538 568146 297774
rect 568382 297538 568466 297774
rect 568702 297538 568734 297774
rect 568114 297454 568734 297538
rect 568114 297218 568146 297454
rect 568382 297218 568466 297454
rect 568702 297218 568734 297454
rect 568114 263774 568734 297218
rect 568114 263538 568146 263774
rect 568382 263538 568466 263774
rect 568702 263538 568734 263774
rect 568114 263454 568734 263538
rect 568114 263218 568146 263454
rect 568382 263218 568466 263454
rect 568702 263218 568734 263454
rect 568114 229774 568734 263218
rect 568114 229538 568146 229774
rect 568382 229538 568466 229774
rect 568702 229538 568734 229774
rect 568114 229454 568734 229538
rect 568114 229218 568146 229454
rect 568382 229218 568466 229454
rect 568702 229218 568734 229454
rect 568114 195774 568734 229218
rect 568114 195538 568146 195774
rect 568382 195538 568466 195774
rect 568702 195538 568734 195774
rect 568114 195454 568734 195538
rect 568114 195218 568146 195454
rect 568382 195218 568466 195454
rect 568702 195218 568734 195454
rect 568114 161774 568734 195218
rect 568114 161538 568146 161774
rect 568382 161538 568466 161774
rect 568702 161538 568734 161774
rect 568114 161454 568734 161538
rect 568114 161218 568146 161454
rect 568382 161218 568466 161454
rect 568702 161218 568734 161454
rect 568114 127774 568734 161218
rect 568114 127538 568146 127774
rect 568382 127538 568466 127774
rect 568702 127538 568734 127774
rect 568114 127454 568734 127538
rect 568114 127218 568146 127454
rect 568382 127218 568466 127454
rect 568702 127218 568734 127454
rect 568114 93774 568734 127218
rect 568114 93538 568146 93774
rect 568382 93538 568466 93774
rect 568702 93538 568734 93774
rect 568114 93454 568734 93538
rect 568114 93218 568146 93454
rect 568382 93218 568466 93454
rect 568702 93218 568734 93454
rect 568114 59774 568734 93218
rect 568114 59538 568146 59774
rect 568382 59538 568466 59774
rect 568702 59538 568734 59774
rect 568114 59454 568734 59538
rect 568114 59218 568146 59454
rect 568382 59218 568466 59454
rect 568702 59218 568734 59454
rect 568114 25774 568734 59218
rect 568114 25538 568146 25774
rect 568382 25538 568466 25774
rect 568702 25538 568734 25774
rect 568114 25454 568734 25538
rect 568114 25218 568146 25454
rect 568382 25218 568466 25454
rect 568702 25218 568734 25454
rect 568114 -6106 568734 25218
rect 568114 -6342 568146 -6106
rect 568382 -6342 568466 -6106
rect 568702 -6342 568734 -6106
rect 568114 -6426 568734 -6342
rect 568114 -6662 568146 -6426
rect 568382 -6662 568466 -6426
rect 568702 -6662 568734 -6426
rect 568114 -7654 568734 -6662
rect 571834 711558 572454 711590
rect 571834 711322 571866 711558
rect 572102 711322 572186 711558
rect 572422 711322 572454 711558
rect 571834 711238 572454 711322
rect 571834 711002 571866 711238
rect 572102 711002 572186 711238
rect 572422 711002 572454 711238
rect 571834 675494 572454 711002
rect 571834 675258 571866 675494
rect 572102 675258 572186 675494
rect 572422 675258 572454 675494
rect 571834 675174 572454 675258
rect 571834 674938 571866 675174
rect 572102 674938 572186 675174
rect 572422 674938 572454 675174
rect 571834 641494 572454 674938
rect 571834 641258 571866 641494
rect 572102 641258 572186 641494
rect 572422 641258 572454 641494
rect 571834 641174 572454 641258
rect 571834 640938 571866 641174
rect 572102 640938 572186 641174
rect 572422 640938 572454 641174
rect 571834 607494 572454 640938
rect 571834 607258 571866 607494
rect 572102 607258 572186 607494
rect 572422 607258 572454 607494
rect 571834 607174 572454 607258
rect 571834 606938 571866 607174
rect 572102 606938 572186 607174
rect 572422 606938 572454 607174
rect 571834 573494 572454 606938
rect 571834 573258 571866 573494
rect 572102 573258 572186 573494
rect 572422 573258 572454 573494
rect 571834 573174 572454 573258
rect 571834 572938 571866 573174
rect 572102 572938 572186 573174
rect 572422 572938 572454 573174
rect 571834 539494 572454 572938
rect 571834 539258 571866 539494
rect 572102 539258 572186 539494
rect 572422 539258 572454 539494
rect 571834 539174 572454 539258
rect 571834 538938 571866 539174
rect 572102 538938 572186 539174
rect 572422 538938 572454 539174
rect 571834 505494 572454 538938
rect 571834 505258 571866 505494
rect 572102 505258 572186 505494
rect 572422 505258 572454 505494
rect 571834 505174 572454 505258
rect 571834 504938 571866 505174
rect 572102 504938 572186 505174
rect 572422 504938 572454 505174
rect 571834 471494 572454 504938
rect 571834 471258 571866 471494
rect 572102 471258 572186 471494
rect 572422 471258 572454 471494
rect 571834 471174 572454 471258
rect 571834 470938 571866 471174
rect 572102 470938 572186 471174
rect 572422 470938 572454 471174
rect 571834 437494 572454 470938
rect 571834 437258 571866 437494
rect 572102 437258 572186 437494
rect 572422 437258 572454 437494
rect 571834 437174 572454 437258
rect 571834 436938 571866 437174
rect 572102 436938 572186 437174
rect 572422 436938 572454 437174
rect 571834 403494 572454 436938
rect 571834 403258 571866 403494
rect 572102 403258 572186 403494
rect 572422 403258 572454 403494
rect 571834 403174 572454 403258
rect 571834 402938 571866 403174
rect 572102 402938 572186 403174
rect 572422 402938 572454 403174
rect 571834 369494 572454 402938
rect 571834 369258 571866 369494
rect 572102 369258 572186 369494
rect 572422 369258 572454 369494
rect 571834 369174 572454 369258
rect 571834 368938 571866 369174
rect 572102 368938 572186 369174
rect 572422 368938 572454 369174
rect 571834 335494 572454 368938
rect 571834 335258 571866 335494
rect 572102 335258 572186 335494
rect 572422 335258 572454 335494
rect 571834 335174 572454 335258
rect 571834 334938 571866 335174
rect 572102 334938 572186 335174
rect 572422 334938 572454 335174
rect 571834 301494 572454 334938
rect 571834 301258 571866 301494
rect 572102 301258 572186 301494
rect 572422 301258 572454 301494
rect 571834 301174 572454 301258
rect 571834 300938 571866 301174
rect 572102 300938 572186 301174
rect 572422 300938 572454 301174
rect 571834 267494 572454 300938
rect 571834 267258 571866 267494
rect 572102 267258 572186 267494
rect 572422 267258 572454 267494
rect 571834 267174 572454 267258
rect 571834 266938 571866 267174
rect 572102 266938 572186 267174
rect 572422 266938 572454 267174
rect 571834 233494 572454 266938
rect 571834 233258 571866 233494
rect 572102 233258 572186 233494
rect 572422 233258 572454 233494
rect 571834 233174 572454 233258
rect 571834 232938 571866 233174
rect 572102 232938 572186 233174
rect 572422 232938 572454 233174
rect 571834 199494 572454 232938
rect 571834 199258 571866 199494
rect 572102 199258 572186 199494
rect 572422 199258 572454 199494
rect 571834 199174 572454 199258
rect 571834 198938 571866 199174
rect 572102 198938 572186 199174
rect 572422 198938 572454 199174
rect 571834 165494 572454 198938
rect 571834 165258 571866 165494
rect 572102 165258 572186 165494
rect 572422 165258 572454 165494
rect 571834 165174 572454 165258
rect 571834 164938 571866 165174
rect 572102 164938 572186 165174
rect 572422 164938 572454 165174
rect 571834 131494 572454 164938
rect 571834 131258 571866 131494
rect 572102 131258 572186 131494
rect 572422 131258 572454 131494
rect 571834 131174 572454 131258
rect 571834 130938 571866 131174
rect 572102 130938 572186 131174
rect 572422 130938 572454 131174
rect 571834 97494 572454 130938
rect 571834 97258 571866 97494
rect 572102 97258 572186 97494
rect 572422 97258 572454 97494
rect 571834 97174 572454 97258
rect 571834 96938 571866 97174
rect 572102 96938 572186 97174
rect 572422 96938 572454 97174
rect 571834 63494 572454 96938
rect 571834 63258 571866 63494
rect 572102 63258 572186 63494
rect 572422 63258 572454 63494
rect 571834 63174 572454 63258
rect 571834 62938 571866 63174
rect 572102 62938 572186 63174
rect 572422 62938 572454 63174
rect 571834 29494 572454 62938
rect 571834 29258 571866 29494
rect 572102 29258 572186 29494
rect 572422 29258 572454 29494
rect 571834 29174 572454 29258
rect 571834 28938 571866 29174
rect 572102 28938 572186 29174
rect 572422 28938 572454 29174
rect 571834 -7066 572454 28938
rect 571834 -7302 571866 -7066
rect 572102 -7302 572186 -7066
rect 572422 -7302 572454 -7066
rect 571834 -7386 572454 -7302
rect 571834 -7622 571866 -7386
rect 572102 -7622 572186 -7386
rect 572422 -7622 572454 -7386
rect 571834 -7654 572454 -7622
rect 579794 704838 580414 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 579794 704602 579826 704838
rect 580062 704602 580146 704838
rect 580382 704602 580414 704838
rect 579794 704518 580414 704602
rect 579794 704282 579826 704518
rect 580062 704282 580146 704518
rect 580382 704282 580414 704518
rect 579794 683454 580414 704282
rect 579794 683218 579826 683454
rect 580062 683218 580146 683454
rect 580382 683218 580414 683454
rect 579794 683134 580414 683218
rect 579794 682898 579826 683134
rect 580062 682898 580146 683134
rect 580382 682898 580414 683134
rect 579794 649454 580414 682898
rect 579794 649218 579826 649454
rect 580062 649218 580146 649454
rect 580382 649218 580414 649454
rect 579794 649134 580414 649218
rect 579794 648898 579826 649134
rect 580062 648898 580146 649134
rect 580382 648898 580414 649134
rect 579794 615454 580414 648898
rect 579794 615218 579826 615454
rect 580062 615218 580146 615454
rect 580382 615218 580414 615454
rect 579794 615134 580414 615218
rect 579794 614898 579826 615134
rect 580062 614898 580146 615134
rect 580382 614898 580414 615134
rect 579794 581454 580414 614898
rect 579794 581218 579826 581454
rect 580062 581218 580146 581454
rect 580382 581218 580414 581454
rect 579794 581134 580414 581218
rect 579794 580898 579826 581134
rect 580062 580898 580146 581134
rect 580382 580898 580414 581134
rect 579794 547454 580414 580898
rect 579794 547218 579826 547454
rect 580062 547218 580146 547454
rect 580382 547218 580414 547454
rect 579794 547134 580414 547218
rect 579794 546898 579826 547134
rect 580062 546898 580146 547134
rect 580382 546898 580414 547134
rect 579794 513454 580414 546898
rect 579794 513218 579826 513454
rect 580062 513218 580146 513454
rect 580382 513218 580414 513454
rect 579794 513134 580414 513218
rect 579794 512898 579826 513134
rect 580062 512898 580146 513134
rect 580382 512898 580414 513134
rect 579794 479454 580414 512898
rect 579794 479218 579826 479454
rect 580062 479218 580146 479454
rect 580382 479218 580414 479454
rect 579794 479134 580414 479218
rect 579794 478898 579826 479134
rect 580062 478898 580146 479134
rect 580382 478898 580414 479134
rect 579794 445454 580414 478898
rect 579794 445218 579826 445454
rect 580062 445218 580146 445454
rect 580382 445218 580414 445454
rect 579794 445134 580414 445218
rect 579794 444898 579826 445134
rect 580062 444898 580146 445134
rect 580382 444898 580414 445134
rect 579794 411454 580414 444898
rect 579794 411218 579826 411454
rect 580062 411218 580146 411454
rect 580382 411218 580414 411454
rect 579794 411134 580414 411218
rect 579794 410898 579826 411134
rect 580062 410898 580146 411134
rect 580382 410898 580414 411134
rect 579794 377454 580414 410898
rect 579794 377218 579826 377454
rect 580062 377218 580146 377454
rect 580382 377218 580414 377454
rect 579794 377134 580414 377218
rect 579794 376898 579826 377134
rect 580062 376898 580146 377134
rect 580382 376898 580414 377134
rect 579794 343454 580414 376898
rect 579794 343218 579826 343454
rect 580062 343218 580146 343454
rect 580382 343218 580414 343454
rect 579794 343134 580414 343218
rect 579794 342898 579826 343134
rect 580062 342898 580146 343134
rect 580382 342898 580414 343134
rect 579794 309454 580414 342898
rect 579794 309218 579826 309454
rect 580062 309218 580146 309454
rect 580382 309218 580414 309454
rect 579794 309134 580414 309218
rect 579794 308898 579826 309134
rect 580062 308898 580146 309134
rect 580382 308898 580414 309134
rect 579794 275454 580414 308898
rect 579794 275218 579826 275454
rect 580062 275218 580146 275454
rect 580382 275218 580414 275454
rect 579794 275134 580414 275218
rect 579794 274898 579826 275134
rect 580062 274898 580146 275134
rect 580382 274898 580414 275134
rect 579794 241454 580414 274898
rect 579794 241218 579826 241454
rect 580062 241218 580146 241454
rect 580382 241218 580414 241454
rect 579794 241134 580414 241218
rect 579794 240898 579826 241134
rect 580062 240898 580146 241134
rect 580382 240898 580414 241134
rect 579794 207454 580414 240898
rect 579794 207218 579826 207454
rect 580062 207218 580146 207454
rect 580382 207218 580414 207454
rect 579794 207134 580414 207218
rect 579794 206898 579826 207134
rect 580062 206898 580146 207134
rect 580382 206898 580414 207134
rect 579794 173454 580414 206898
rect 579794 173218 579826 173454
rect 580062 173218 580146 173454
rect 580382 173218 580414 173454
rect 579794 173134 580414 173218
rect 579794 172898 579826 173134
rect 580062 172898 580146 173134
rect 580382 172898 580414 173134
rect 579794 139454 580414 172898
rect 579794 139218 579826 139454
rect 580062 139218 580146 139454
rect 580382 139218 580414 139454
rect 579794 139134 580414 139218
rect 579794 138898 579826 139134
rect 580062 138898 580146 139134
rect 580382 138898 580414 139134
rect 579794 105454 580414 138898
rect 579794 105218 579826 105454
rect 580062 105218 580146 105454
rect 580382 105218 580414 105454
rect 579794 105134 580414 105218
rect 579794 104898 579826 105134
rect 580062 104898 580146 105134
rect 580382 104898 580414 105134
rect 579794 71454 580414 104898
rect 579794 71218 579826 71454
rect 580062 71218 580146 71454
rect 580382 71218 580414 71454
rect 579794 71134 580414 71218
rect 579794 70898 579826 71134
rect 580062 70898 580146 71134
rect 580382 70898 580414 71134
rect 579794 37454 580414 70898
rect 579794 37218 579826 37454
rect 580062 37218 580146 37454
rect 580382 37218 580414 37454
rect 579794 37134 580414 37218
rect 579794 36898 579826 37134
rect 580062 36898 580146 37134
rect 580382 36898 580414 37134
rect 579794 3454 580414 36898
rect 579794 3218 579826 3454
rect 580062 3218 580146 3454
rect 580382 3218 580414 3454
rect 579794 3134 580414 3218
rect 579794 2898 579826 3134
rect 580062 2898 580146 3134
rect 580382 2898 580414 3134
rect 579794 -346 580414 2898
rect 579794 -582 579826 -346
rect 580062 -582 580146 -346
rect 580382 -582 580414 -346
rect 579794 -666 580414 -582
rect 579794 -902 579826 -666
rect 580062 -902 580146 -666
rect 580382 -902 580414 -666
rect 579794 -7654 580414 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 683454 585930 704282
rect 585310 683218 585342 683454
rect 585578 683218 585662 683454
rect 585898 683218 585930 683454
rect 585310 683134 585930 683218
rect 585310 682898 585342 683134
rect 585578 682898 585662 683134
rect 585898 682898 585930 683134
rect 585310 649454 585930 682898
rect 585310 649218 585342 649454
rect 585578 649218 585662 649454
rect 585898 649218 585930 649454
rect 585310 649134 585930 649218
rect 585310 648898 585342 649134
rect 585578 648898 585662 649134
rect 585898 648898 585930 649134
rect 585310 615454 585930 648898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 581454 585930 614898
rect 585310 581218 585342 581454
rect 585578 581218 585662 581454
rect 585898 581218 585930 581454
rect 585310 581134 585930 581218
rect 585310 580898 585342 581134
rect 585578 580898 585662 581134
rect 585898 580898 585930 581134
rect 585310 547454 585930 580898
rect 585310 547218 585342 547454
rect 585578 547218 585662 547454
rect 585898 547218 585930 547454
rect 585310 547134 585930 547218
rect 585310 546898 585342 547134
rect 585578 546898 585662 547134
rect 585898 546898 585930 547134
rect 585310 513454 585930 546898
rect 585310 513218 585342 513454
rect 585578 513218 585662 513454
rect 585898 513218 585930 513454
rect 585310 513134 585930 513218
rect 585310 512898 585342 513134
rect 585578 512898 585662 513134
rect 585898 512898 585930 513134
rect 585310 479454 585930 512898
rect 585310 479218 585342 479454
rect 585578 479218 585662 479454
rect 585898 479218 585930 479454
rect 585310 479134 585930 479218
rect 585310 478898 585342 479134
rect 585578 478898 585662 479134
rect 585898 478898 585930 479134
rect 585310 445454 585930 478898
rect 585310 445218 585342 445454
rect 585578 445218 585662 445454
rect 585898 445218 585930 445454
rect 585310 445134 585930 445218
rect 585310 444898 585342 445134
rect 585578 444898 585662 445134
rect 585898 444898 585930 445134
rect 585310 411454 585930 444898
rect 585310 411218 585342 411454
rect 585578 411218 585662 411454
rect 585898 411218 585930 411454
rect 585310 411134 585930 411218
rect 585310 410898 585342 411134
rect 585578 410898 585662 411134
rect 585898 410898 585930 411134
rect 585310 377454 585930 410898
rect 585310 377218 585342 377454
rect 585578 377218 585662 377454
rect 585898 377218 585930 377454
rect 585310 377134 585930 377218
rect 585310 376898 585342 377134
rect 585578 376898 585662 377134
rect 585898 376898 585930 377134
rect 585310 343454 585930 376898
rect 585310 343218 585342 343454
rect 585578 343218 585662 343454
rect 585898 343218 585930 343454
rect 585310 343134 585930 343218
rect 585310 342898 585342 343134
rect 585578 342898 585662 343134
rect 585898 342898 585930 343134
rect 585310 309454 585930 342898
rect 585310 309218 585342 309454
rect 585578 309218 585662 309454
rect 585898 309218 585930 309454
rect 585310 309134 585930 309218
rect 585310 308898 585342 309134
rect 585578 308898 585662 309134
rect 585898 308898 585930 309134
rect 585310 275454 585930 308898
rect 585310 275218 585342 275454
rect 585578 275218 585662 275454
rect 585898 275218 585930 275454
rect 585310 275134 585930 275218
rect 585310 274898 585342 275134
rect 585578 274898 585662 275134
rect 585898 274898 585930 275134
rect 585310 241454 585930 274898
rect 585310 241218 585342 241454
rect 585578 241218 585662 241454
rect 585898 241218 585930 241454
rect 585310 241134 585930 241218
rect 585310 240898 585342 241134
rect 585578 240898 585662 241134
rect 585898 240898 585930 241134
rect 585310 207454 585930 240898
rect 585310 207218 585342 207454
rect 585578 207218 585662 207454
rect 585898 207218 585930 207454
rect 585310 207134 585930 207218
rect 585310 206898 585342 207134
rect 585578 206898 585662 207134
rect 585898 206898 585930 207134
rect 585310 173454 585930 206898
rect 585310 173218 585342 173454
rect 585578 173218 585662 173454
rect 585898 173218 585930 173454
rect 585310 173134 585930 173218
rect 585310 172898 585342 173134
rect 585578 172898 585662 173134
rect 585898 172898 585930 173134
rect 585310 139454 585930 172898
rect 585310 139218 585342 139454
rect 585578 139218 585662 139454
rect 585898 139218 585930 139454
rect 585310 139134 585930 139218
rect 585310 138898 585342 139134
rect 585578 138898 585662 139134
rect 585898 138898 585930 139134
rect 585310 105454 585930 138898
rect 585310 105218 585342 105454
rect 585578 105218 585662 105454
rect 585898 105218 585930 105454
rect 585310 105134 585930 105218
rect 585310 104898 585342 105134
rect 585578 104898 585662 105134
rect 585898 104898 585930 105134
rect 585310 71454 585930 104898
rect 585310 71218 585342 71454
rect 585578 71218 585662 71454
rect 585898 71218 585930 71454
rect 585310 71134 585930 71218
rect 585310 70898 585342 71134
rect 585578 70898 585662 71134
rect 585898 70898 585930 71134
rect 585310 37454 585930 70898
rect 585310 37218 585342 37454
rect 585578 37218 585662 37454
rect 585898 37218 585930 37454
rect 585310 37134 585930 37218
rect 585310 36898 585342 37134
rect 585578 36898 585662 37134
rect 585898 36898 585930 37134
rect 585310 3454 585930 36898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 687174 586890 705242
rect 586270 686938 586302 687174
rect 586538 686938 586622 687174
rect 586858 686938 586890 687174
rect 586270 686854 586890 686938
rect 586270 686618 586302 686854
rect 586538 686618 586622 686854
rect 586858 686618 586890 686854
rect 586270 653174 586890 686618
rect 586270 652938 586302 653174
rect 586538 652938 586622 653174
rect 586858 652938 586890 653174
rect 586270 652854 586890 652938
rect 586270 652618 586302 652854
rect 586538 652618 586622 652854
rect 586858 652618 586890 652854
rect 586270 619174 586890 652618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 585174 586890 618618
rect 586270 584938 586302 585174
rect 586538 584938 586622 585174
rect 586858 584938 586890 585174
rect 586270 584854 586890 584938
rect 586270 584618 586302 584854
rect 586538 584618 586622 584854
rect 586858 584618 586890 584854
rect 586270 551174 586890 584618
rect 586270 550938 586302 551174
rect 586538 550938 586622 551174
rect 586858 550938 586890 551174
rect 586270 550854 586890 550938
rect 586270 550618 586302 550854
rect 586538 550618 586622 550854
rect 586858 550618 586890 550854
rect 586270 517174 586890 550618
rect 586270 516938 586302 517174
rect 586538 516938 586622 517174
rect 586858 516938 586890 517174
rect 586270 516854 586890 516938
rect 586270 516618 586302 516854
rect 586538 516618 586622 516854
rect 586858 516618 586890 516854
rect 586270 483174 586890 516618
rect 586270 482938 586302 483174
rect 586538 482938 586622 483174
rect 586858 482938 586890 483174
rect 586270 482854 586890 482938
rect 586270 482618 586302 482854
rect 586538 482618 586622 482854
rect 586858 482618 586890 482854
rect 586270 449174 586890 482618
rect 586270 448938 586302 449174
rect 586538 448938 586622 449174
rect 586858 448938 586890 449174
rect 586270 448854 586890 448938
rect 586270 448618 586302 448854
rect 586538 448618 586622 448854
rect 586858 448618 586890 448854
rect 586270 415174 586890 448618
rect 586270 414938 586302 415174
rect 586538 414938 586622 415174
rect 586858 414938 586890 415174
rect 586270 414854 586890 414938
rect 586270 414618 586302 414854
rect 586538 414618 586622 414854
rect 586858 414618 586890 414854
rect 586270 381174 586890 414618
rect 586270 380938 586302 381174
rect 586538 380938 586622 381174
rect 586858 380938 586890 381174
rect 586270 380854 586890 380938
rect 586270 380618 586302 380854
rect 586538 380618 586622 380854
rect 586858 380618 586890 380854
rect 586270 347174 586890 380618
rect 586270 346938 586302 347174
rect 586538 346938 586622 347174
rect 586858 346938 586890 347174
rect 586270 346854 586890 346938
rect 586270 346618 586302 346854
rect 586538 346618 586622 346854
rect 586858 346618 586890 346854
rect 586270 313174 586890 346618
rect 586270 312938 586302 313174
rect 586538 312938 586622 313174
rect 586858 312938 586890 313174
rect 586270 312854 586890 312938
rect 586270 312618 586302 312854
rect 586538 312618 586622 312854
rect 586858 312618 586890 312854
rect 586270 279174 586890 312618
rect 586270 278938 586302 279174
rect 586538 278938 586622 279174
rect 586858 278938 586890 279174
rect 586270 278854 586890 278938
rect 586270 278618 586302 278854
rect 586538 278618 586622 278854
rect 586858 278618 586890 278854
rect 586270 245174 586890 278618
rect 586270 244938 586302 245174
rect 586538 244938 586622 245174
rect 586858 244938 586890 245174
rect 586270 244854 586890 244938
rect 586270 244618 586302 244854
rect 586538 244618 586622 244854
rect 586858 244618 586890 244854
rect 586270 211174 586890 244618
rect 586270 210938 586302 211174
rect 586538 210938 586622 211174
rect 586858 210938 586890 211174
rect 586270 210854 586890 210938
rect 586270 210618 586302 210854
rect 586538 210618 586622 210854
rect 586858 210618 586890 210854
rect 586270 177174 586890 210618
rect 586270 176938 586302 177174
rect 586538 176938 586622 177174
rect 586858 176938 586890 177174
rect 586270 176854 586890 176938
rect 586270 176618 586302 176854
rect 586538 176618 586622 176854
rect 586858 176618 586890 176854
rect 586270 143174 586890 176618
rect 586270 142938 586302 143174
rect 586538 142938 586622 143174
rect 586858 142938 586890 143174
rect 586270 142854 586890 142938
rect 586270 142618 586302 142854
rect 586538 142618 586622 142854
rect 586858 142618 586890 142854
rect 586270 109174 586890 142618
rect 586270 108938 586302 109174
rect 586538 108938 586622 109174
rect 586858 108938 586890 109174
rect 586270 108854 586890 108938
rect 586270 108618 586302 108854
rect 586538 108618 586622 108854
rect 586858 108618 586890 108854
rect 586270 75174 586890 108618
rect 586270 74938 586302 75174
rect 586538 74938 586622 75174
rect 586858 74938 586890 75174
rect 586270 74854 586890 74938
rect 586270 74618 586302 74854
rect 586538 74618 586622 74854
rect 586858 74618 586890 74854
rect 586270 41174 586890 74618
rect 586270 40938 586302 41174
rect 586538 40938 586622 41174
rect 586858 40938 586890 41174
rect 586270 40854 586890 40938
rect 586270 40618 586302 40854
rect 586538 40618 586622 40854
rect 586858 40618 586890 40854
rect 586270 7174 586890 40618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 690894 587850 706202
rect 587230 690658 587262 690894
rect 587498 690658 587582 690894
rect 587818 690658 587850 690894
rect 587230 690574 587850 690658
rect 587230 690338 587262 690574
rect 587498 690338 587582 690574
rect 587818 690338 587850 690574
rect 587230 656894 587850 690338
rect 587230 656658 587262 656894
rect 587498 656658 587582 656894
rect 587818 656658 587850 656894
rect 587230 656574 587850 656658
rect 587230 656338 587262 656574
rect 587498 656338 587582 656574
rect 587818 656338 587850 656574
rect 587230 622894 587850 656338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 588894 587850 622338
rect 587230 588658 587262 588894
rect 587498 588658 587582 588894
rect 587818 588658 587850 588894
rect 587230 588574 587850 588658
rect 587230 588338 587262 588574
rect 587498 588338 587582 588574
rect 587818 588338 587850 588574
rect 587230 554894 587850 588338
rect 587230 554658 587262 554894
rect 587498 554658 587582 554894
rect 587818 554658 587850 554894
rect 587230 554574 587850 554658
rect 587230 554338 587262 554574
rect 587498 554338 587582 554574
rect 587818 554338 587850 554574
rect 587230 520894 587850 554338
rect 587230 520658 587262 520894
rect 587498 520658 587582 520894
rect 587818 520658 587850 520894
rect 587230 520574 587850 520658
rect 587230 520338 587262 520574
rect 587498 520338 587582 520574
rect 587818 520338 587850 520574
rect 587230 486894 587850 520338
rect 587230 486658 587262 486894
rect 587498 486658 587582 486894
rect 587818 486658 587850 486894
rect 587230 486574 587850 486658
rect 587230 486338 587262 486574
rect 587498 486338 587582 486574
rect 587818 486338 587850 486574
rect 587230 452894 587850 486338
rect 587230 452658 587262 452894
rect 587498 452658 587582 452894
rect 587818 452658 587850 452894
rect 587230 452574 587850 452658
rect 587230 452338 587262 452574
rect 587498 452338 587582 452574
rect 587818 452338 587850 452574
rect 587230 418894 587850 452338
rect 587230 418658 587262 418894
rect 587498 418658 587582 418894
rect 587818 418658 587850 418894
rect 587230 418574 587850 418658
rect 587230 418338 587262 418574
rect 587498 418338 587582 418574
rect 587818 418338 587850 418574
rect 587230 384894 587850 418338
rect 587230 384658 587262 384894
rect 587498 384658 587582 384894
rect 587818 384658 587850 384894
rect 587230 384574 587850 384658
rect 587230 384338 587262 384574
rect 587498 384338 587582 384574
rect 587818 384338 587850 384574
rect 587230 350894 587850 384338
rect 587230 350658 587262 350894
rect 587498 350658 587582 350894
rect 587818 350658 587850 350894
rect 587230 350574 587850 350658
rect 587230 350338 587262 350574
rect 587498 350338 587582 350574
rect 587818 350338 587850 350574
rect 587230 316894 587850 350338
rect 587230 316658 587262 316894
rect 587498 316658 587582 316894
rect 587818 316658 587850 316894
rect 587230 316574 587850 316658
rect 587230 316338 587262 316574
rect 587498 316338 587582 316574
rect 587818 316338 587850 316574
rect 587230 282894 587850 316338
rect 587230 282658 587262 282894
rect 587498 282658 587582 282894
rect 587818 282658 587850 282894
rect 587230 282574 587850 282658
rect 587230 282338 587262 282574
rect 587498 282338 587582 282574
rect 587818 282338 587850 282574
rect 587230 248894 587850 282338
rect 587230 248658 587262 248894
rect 587498 248658 587582 248894
rect 587818 248658 587850 248894
rect 587230 248574 587850 248658
rect 587230 248338 587262 248574
rect 587498 248338 587582 248574
rect 587818 248338 587850 248574
rect 587230 214894 587850 248338
rect 587230 214658 587262 214894
rect 587498 214658 587582 214894
rect 587818 214658 587850 214894
rect 587230 214574 587850 214658
rect 587230 214338 587262 214574
rect 587498 214338 587582 214574
rect 587818 214338 587850 214574
rect 587230 180894 587850 214338
rect 587230 180658 587262 180894
rect 587498 180658 587582 180894
rect 587818 180658 587850 180894
rect 587230 180574 587850 180658
rect 587230 180338 587262 180574
rect 587498 180338 587582 180574
rect 587818 180338 587850 180574
rect 587230 146894 587850 180338
rect 587230 146658 587262 146894
rect 587498 146658 587582 146894
rect 587818 146658 587850 146894
rect 587230 146574 587850 146658
rect 587230 146338 587262 146574
rect 587498 146338 587582 146574
rect 587818 146338 587850 146574
rect 587230 112894 587850 146338
rect 587230 112658 587262 112894
rect 587498 112658 587582 112894
rect 587818 112658 587850 112894
rect 587230 112574 587850 112658
rect 587230 112338 587262 112574
rect 587498 112338 587582 112574
rect 587818 112338 587850 112574
rect 587230 78894 587850 112338
rect 587230 78658 587262 78894
rect 587498 78658 587582 78894
rect 587818 78658 587850 78894
rect 587230 78574 587850 78658
rect 587230 78338 587262 78574
rect 587498 78338 587582 78574
rect 587818 78338 587850 78574
rect 587230 44894 587850 78338
rect 587230 44658 587262 44894
rect 587498 44658 587582 44894
rect 587818 44658 587850 44894
rect 587230 44574 587850 44658
rect 587230 44338 587262 44574
rect 587498 44338 587582 44574
rect 587818 44338 587850 44574
rect 587230 10894 587850 44338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 694614 588810 707162
rect 588190 694378 588222 694614
rect 588458 694378 588542 694614
rect 588778 694378 588810 694614
rect 588190 694294 588810 694378
rect 588190 694058 588222 694294
rect 588458 694058 588542 694294
rect 588778 694058 588810 694294
rect 588190 660614 588810 694058
rect 588190 660378 588222 660614
rect 588458 660378 588542 660614
rect 588778 660378 588810 660614
rect 588190 660294 588810 660378
rect 588190 660058 588222 660294
rect 588458 660058 588542 660294
rect 588778 660058 588810 660294
rect 588190 626614 588810 660058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 592614 588810 626058
rect 588190 592378 588222 592614
rect 588458 592378 588542 592614
rect 588778 592378 588810 592614
rect 588190 592294 588810 592378
rect 588190 592058 588222 592294
rect 588458 592058 588542 592294
rect 588778 592058 588810 592294
rect 588190 558614 588810 592058
rect 588190 558378 588222 558614
rect 588458 558378 588542 558614
rect 588778 558378 588810 558614
rect 588190 558294 588810 558378
rect 588190 558058 588222 558294
rect 588458 558058 588542 558294
rect 588778 558058 588810 558294
rect 588190 524614 588810 558058
rect 588190 524378 588222 524614
rect 588458 524378 588542 524614
rect 588778 524378 588810 524614
rect 588190 524294 588810 524378
rect 588190 524058 588222 524294
rect 588458 524058 588542 524294
rect 588778 524058 588810 524294
rect 588190 490614 588810 524058
rect 588190 490378 588222 490614
rect 588458 490378 588542 490614
rect 588778 490378 588810 490614
rect 588190 490294 588810 490378
rect 588190 490058 588222 490294
rect 588458 490058 588542 490294
rect 588778 490058 588810 490294
rect 588190 456614 588810 490058
rect 588190 456378 588222 456614
rect 588458 456378 588542 456614
rect 588778 456378 588810 456614
rect 588190 456294 588810 456378
rect 588190 456058 588222 456294
rect 588458 456058 588542 456294
rect 588778 456058 588810 456294
rect 588190 422614 588810 456058
rect 588190 422378 588222 422614
rect 588458 422378 588542 422614
rect 588778 422378 588810 422614
rect 588190 422294 588810 422378
rect 588190 422058 588222 422294
rect 588458 422058 588542 422294
rect 588778 422058 588810 422294
rect 588190 388614 588810 422058
rect 588190 388378 588222 388614
rect 588458 388378 588542 388614
rect 588778 388378 588810 388614
rect 588190 388294 588810 388378
rect 588190 388058 588222 388294
rect 588458 388058 588542 388294
rect 588778 388058 588810 388294
rect 588190 354614 588810 388058
rect 588190 354378 588222 354614
rect 588458 354378 588542 354614
rect 588778 354378 588810 354614
rect 588190 354294 588810 354378
rect 588190 354058 588222 354294
rect 588458 354058 588542 354294
rect 588778 354058 588810 354294
rect 588190 320614 588810 354058
rect 588190 320378 588222 320614
rect 588458 320378 588542 320614
rect 588778 320378 588810 320614
rect 588190 320294 588810 320378
rect 588190 320058 588222 320294
rect 588458 320058 588542 320294
rect 588778 320058 588810 320294
rect 588190 286614 588810 320058
rect 588190 286378 588222 286614
rect 588458 286378 588542 286614
rect 588778 286378 588810 286614
rect 588190 286294 588810 286378
rect 588190 286058 588222 286294
rect 588458 286058 588542 286294
rect 588778 286058 588810 286294
rect 588190 252614 588810 286058
rect 588190 252378 588222 252614
rect 588458 252378 588542 252614
rect 588778 252378 588810 252614
rect 588190 252294 588810 252378
rect 588190 252058 588222 252294
rect 588458 252058 588542 252294
rect 588778 252058 588810 252294
rect 588190 218614 588810 252058
rect 588190 218378 588222 218614
rect 588458 218378 588542 218614
rect 588778 218378 588810 218614
rect 588190 218294 588810 218378
rect 588190 218058 588222 218294
rect 588458 218058 588542 218294
rect 588778 218058 588810 218294
rect 588190 184614 588810 218058
rect 588190 184378 588222 184614
rect 588458 184378 588542 184614
rect 588778 184378 588810 184614
rect 588190 184294 588810 184378
rect 588190 184058 588222 184294
rect 588458 184058 588542 184294
rect 588778 184058 588810 184294
rect 588190 150614 588810 184058
rect 588190 150378 588222 150614
rect 588458 150378 588542 150614
rect 588778 150378 588810 150614
rect 588190 150294 588810 150378
rect 588190 150058 588222 150294
rect 588458 150058 588542 150294
rect 588778 150058 588810 150294
rect 588190 116614 588810 150058
rect 588190 116378 588222 116614
rect 588458 116378 588542 116614
rect 588778 116378 588810 116614
rect 588190 116294 588810 116378
rect 588190 116058 588222 116294
rect 588458 116058 588542 116294
rect 588778 116058 588810 116294
rect 588190 82614 588810 116058
rect 588190 82378 588222 82614
rect 588458 82378 588542 82614
rect 588778 82378 588810 82614
rect 588190 82294 588810 82378
rect 588190 82058 588222 82294
rect 588458 82058 588542 82294
rect 588778 82058 588810 82294
rect 588190 48614 588810 82058
rect 588190 48378 588222 48614
rect 588458 48378 588542 48614
rect 588778 48378 588810 48614
rect 588190 48294 588810 48378
rect 588190 48058 588222 48294
rect 588458 48058 588542 48294
rect 588778 48058 588810 48294
rect 588190 14614 588810 48058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 698334 589770 708122
rect 589150 698098 589182 698334
rect 589418 698098 589502 698334
rect 589738 698098 589770 698334
rect 589150 698014 589770 698098
rect 589150 697778 589182 698014
rect 589418 697778 589502 698014
rect 589738 697778 589770 698014
rect 589150 664334 589770 697778
rect 589150 664098 589182 664334
rect 589418 664098 589502 664334
rect 589738 664098 589770 664334
rect 589150 664014 589770 664098
rect 589150 663778 589182 664014
rect 589418 663778 589502 664014
rect 589738 663778 589770 664014
rect 589150 630334 589770 663778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 596334 589770 629778
rect 589150 596098 589182 596334
rect 589418 596098 589502 596334
rect 589738 596098 589770 596334
rect 589150 596014 589770 596098
rect 589150 595778 589182 596014
rect 589418 595778 589502 596014
rect 589738 595778 589770 596014
rect 589150 562334 589770 595778
rect 589150 562098 589182 562334
rect 589418 562098 589502 562334
rect 589738 562098 589770 562334
rect 589150 562014 589770 562098
rect 589150 561778 589182 562014
rect 589418 561778 589502 562014
rect 589738 561778 589770 562014
rect 589150 528334 589770 561778
rect 589150 528098 589182 528334
rect 589418 528098 589502 528334
rect 589738 528098 589770 528334
rect 589150 528014 589770 528098
rect 589150 527778 589182 528014
rect 589418 527778 589502 528014
rect 589738 527778 589770 528014
rect 589150 494334 589770 527778
rect 589150 494098 589182 494334
rect 589418 494098 589502 494334
rect 589738 494098 589770 494334
rect 589150 494014 589770 494098
rect 589150 493778 589182 494014
rect 589418 493778 589502 494014
rect 589738 493778 589770 494014
rect 589150 460334 589770 493778
rect 589150 460098 589182 460334
rect 589418 460098 589502 460334
rect 589738 460098 589770 460334
rect 589150 460014 589770 460098
rect 589150 459778 589182 460014
rect 589418 459778 589502 460014
rect 589738 459778 589770 460014
rect 589150 426334 589770 459778
rect 589150 426098 589182 426334
rect 589418 426098 589502 426334
rect 589738 426098 589770 426334
rect 589150 426014 589770 426098
rect 589150 425778 589182 426014
rect 589418 425778 589502 426014
rect 589738 425778 589770 426014
rect 589150 392334 589770 425778
rect 589150 392098 589182 392334
rect 589418 392098 589502 392334
rect 589738 392098 589770 392334
rect 589150 392014 589770 392098
rect 589150 391778 589182 392014
rect 589418 391778 589502 392014
rect 589738 391778 589770 392014
rect 589150 358334 589770 391778
rect 589150 358098 589182 358334
rect 589418 358098 589502 358334
rect 589738 358098 589770 358334
rect 589150 358014 589770 358098
rect 589150 357778 589182 358014
rect 589418 357778 589502 358014
rect 589738 357778 589770 358014
rect 589150 324334 589770 357778
rect 589150 324098 589182 324334
rect 589418 324098 589502 324334
rect 589738 324098 589770 324334
rect 589150 324014 589770 324098
rect 589150 323778 589182 324014
rect 589418 323778 589502 324014
rect 589738 323778 589770 324014
rect 589150 290334 589770 323778
rect 589150 290098 589182 290334
rect 589418 290098 589502 290334
rect 589738 290098 589770 290334
rect 589150 290014 589770 290098
rect 589150 289778 589182 290014
rect 589418 289778 589502 290014
rect 589738 289778 589770 290014
rect 589150 256334 589770 289778
rect 589150 256098 589182 256334
rect 589418 256098 589502 256334
rect 589738 256098 589770 256334
rect 589150 256014 589770 256098
rect 589150 255778 589182 256014
rect 589418 255778 589502 256014
rect 589738 255778 589770 256014
rect 589150 222334 589770 255778
rect 589150 222098 589182 222334
rect 589418 222098 589502 222334
rect 589738 222098 589770 222334
rect 589150 222014 589770 222098
rect 589150 221778 589182 222014
rect 589418 221778 589502 222014
rect 589738 221778 589770 222014
rect 589150 188334 589770 221778
rect 589150 188098 589182 188334
rect 589418 188098 589502 188334
rect 589738 188098 589770 188334
rect 589150 188014 589770 188098
rect 589150 187778 589182 188014
rect 589418 187778 589502 188014
rect 589738 187778 589770 188014
rect 589150 154334 589770 187778
rect 589150 154098 589182 154334
rect 589418 154098 589502 154334
rect 589738 154098 589770 154334
rect 589150 154014 589770 154098
rect 589150 153778 589182 154014
rect 589418 153778 589502 154014
rect 589738 153778 589770 154014
rect 589150 120334 589770 153778
rect 589150 120098 589182 120334
rect 589418 120098 589502 120334
rect 589738 120098 589770 120334
rect 589150 120014 589770 120098
rect 589150 119778 589182 120014
rect 589418 119778 589502 120014
rect 589738 119778 589770 120014
rect 589150 86334 589770 119778
rect 589150 86098 589182 86334
rect 589418 86098 589502 86334
rect 589738 86098 589770 86334
rect 589150 86014 589770 86098
rect 589150 85778 589182 86014
rect 589418 85778 589502 86014
rect 589738 85778 589770 86014
rect 589150 52334 589770 85778
rect 589150 52098 589182 52334
rect 589418 52098 589502 52334
rect 589738 52098 589770 52334
rect 589150 52014 589770 52098
rect 589150 51778 589182 52014
rect 589418 51778 589502 52014
rect 589738 51778 589770 52014
rect 589150 18334 589770 51778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 668054 590730 709082
rect 590110 667818 590142 668054
rect 590378 667818 590462 668054
rect 590698 667818 590730 668054
rect 590110 667734 590730 667818
rect 590110 667498 590142 667734
rect 590378 667498 590462 667734
rect 590698 667498 590730 667734
rect 590110 634054 590730 667498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 600054 590730 633498
rect 590110 599818 590142 600054
rect 590378 599818 590462 600054
rect 590698 599818 590730 600054
rect 590110 599734 590730 599818
rect 590110 599498 590142 599734
rect 590378 599498 590462 599734
rect 590698 599498 590730 599734
rect 590110 566054 590730 599498
rect 590110 565818 590142 566054
rect 590378 565818 590462 566054
rect 590698 565818 590730 566054
rect 590110 565734 590730 565818
rect 590110 565498 590142 565734
rect 590378 565498 590462 565734
rect 590698 565498 590730 565734
rect 590110 532054 590730 565498
rect 590110 531818 590142 532054
rect 590378 531818 590462 532054
rect 590698 531818 590730 532054
rect 590110 531734 590730 531818
rect 590110 531498 590142 531734
rect 590378 531498 590462 531734
rect 590698 531498 590730 531734
rect 590110 498054 590730 531498
rect 590110 497818 590142 498054
rect 590378 497818 590462 498054
rect 590698 497818 590730 498054
rect 590110 497734 590730 497818
rect 590110 497498 590142 497734
rect 590378 497498 590462 497734
rect 590698 497498 590730 497734
rect 590110 464054 590730 497498
rect 590110 463818 590142 464054
rect 590378 463818 590462 464054
rect 590698 463818 590730 464054
rect 590110 463734 590730 463818
rect 590110 463498 590142 463734
rect 590378 463498 590462 463734
rect 590698 463498 590730 463734
rect 590110 430054 590730 463498
rect 590110 429818 590142 430054
rect 590378 429818 590462 430054
rect 590698 429818 590730 430054
rect 590110 429734 590730 429818
rect 590110 429498 590142 429734
rect 590378 429498 590462 429734
rect 590698 429498 590730 429734
rect 590110 396054 590730 429498
rect 590110 395818 590142 396054
rect 590378 395818 590462 396054
rect 590698 395818 590730 396054
rect 590110 395734 590730 395818
rect 590110 395498 590142 395734
rect 590378 395498 590462 395734
rect 590698 395498 590730 395734
rect 590110 362054 590730 395498
rect 590110 361818 590142 362054
rect 590378 361818 590462 362054
rect 590698 361818 590730 362054
rect 590110 361734 590730 361818
rect 590110 361498 590142 361734
rect 590378 361498 590462 361734
rect 590698 361498 590730 361734
rect 590110 328054 590730 361498
rect 590110 327818 590142 328054
rect 590378 327818 590462 328054
rect 590698 327818 590730 328054
rect 590110 327734 590730 327818
rect 590110 327498 590142 327734
rect 590378 327498 590462 327734
rect 590698 327498 590730 327734
rect 590110 294054 590730 327498
rect 590110 293818 590142 294054
rect 590378 293818 590462 294054
rect 590698 293818 590730 294054
rect 590110 293734 590730 293818
rect 590110 293498 590142 293734
rect 590378 293498 590462 293734
rect 590698 293498 590730 293734
rect 590110 260054 590730 293498
rect 590110 259818 590142 260054
rect 590378 259818 590462 260054
rect 590698 259818 590730 260054
rect 590110 259734 590730 259818
rect 590110 259498 590142 259734
rect 590378 259498 590462 259734
rect 590698 259498 590730 259734
rect 590110 226054 590730 259498
rect 590110 225818 590142 226054
rect 590378 225818 590462 226054
rect 590698 225818 590730 226054
rect 590110 225734 590730 225818
rect 590110 225498 590142 225734
rect 590378 225498 590462 225734
rect 590698 225498 590730 225734
rect 590110 192054 590730 225498
rect 590110 191818 590142 192054
rect 590378 191818 590462 192054
rect 590698 191818 590730 192054
rect 590110 191734 590730 191818
rect 590110 191498 590142 191734
rect 590378 191498 590462 191734
rect 590698 191498 590730 191734
rect 590110 158054 590730 191498
rect 590110 157818 590142 158054
rect 590378 157818 590462 158054
rect 590698 157818 590730 158054
rect 590110 157734 590730 157818
rect 590110 157498 590142 157734
rect 590378 157498 590462 157734
rect 590698 157498 590730 157734
rect 590110 124054 590730 157498
rect 590110 123818 590142 124054
rect 590378 123818 590462 124054
rect 590698 123818 590730 124054
rect 590110 123734 590730 123818
rect 590110 123498 590142 123734
rect 590378 123498 590462 123734
rect 590698 123498 590730 123734
rect 590110 90054 590730 123498
rect 590110 89818 590142 90054
rect 590378 89818 590462 90054
rect 590698 89818 590730 90054
rect 590110 89734 590730 89818
rect 590110 89498 590142 89734
rect 590378 89498 590462 89734
rect 590698 89498 590730 89734
rect 590110 56054 590730 89498
rect 590110 55818 590142 56054
rect 590378 55818 590462 56054
rect 590698 55818 590730 56054
rect 590110 55734 590730 55818
rect 590110 55498 590142 55734
rect 590378 55498 590462 55734
rect 590698 55498 590730 55734
rect 590110 22054 590730 55498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 671774 591690 710042
rect 591070 671538 591102 671774
rect 591338 671538 591422 671774
rect 591658 671538 591690 671774
rect 591070 671454 591690 671538
rect 591070 671218 591102 671454
rect 591338 671218 591422 671454
rect 591658 671218 591690 671454
rect 591070 637774 591690 671218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 603774 591690 637218
rect 591070 603538 591102 603774
rect 591338 603538 591422 603774
rect 591658 603538 591690 603774
rect 591070 603454 591690 603538
rect 591070 603218 591102 603454
rect 591338 603218 591422 603454
rect 591658 603218 591690 603454
rect 591070 569774 591690 603218
rect 591070 569538 591102 569774
rect 591338 569538 591422 569774
rect 591658 569538 591690 569774
rect 591070 569454 591690 569538
rect 591070 569218 591102 569454
rect 591338 569218 591422 569454
rect 591658 569218 591690 569454
rect 591070 535774 591690 569218
rect 591070 535538 591102 535774
rect 591338 535538 591422 535774
rect 591658 535538 591690 535774
rect 591070 535454 591690 535538
rect 591070 535218 591102 535454
rect 591338 535218 591422 535454
rect 591658 535218 591690 535454
rect 591070 501774 591690 535218
rect 591070 501538 591102 501774
rect 591338 501538 591422 501774
rect 591658 501538 591690 501774
rect 591070 501454 591690 501538
rect 591070 501218 591102 501454
rect 591338 501218 591422 501454
rect 591658 501218 591690 501454
rect 591070 467774 591690 501218
rect 591070 467538 591102 467774
rect 591338 467538 591422 467774
rect 591658 467538 591690 467774
rect 591070 467454 591690 467538
rect 591070 467218 591102 467454
rect 591338 467218 591422 467454
rect 591658 467218 591690 467454
rect 591070 433774 591690 467218
rect 591070 433538 591102 433774
rect 591338 433538 591422 433774
rect 591658 433538 591690 433774
rect 591070 433454 591690 433538
rect 591070 433218 591102 433454
rect 591338 433218 591422 433454
rect 591658 433218 591690 433454
rect 591070 399774 591690 433218
rect 591070 399538 591102 399774
rect 591338 399538 591422 399774
rect 591658 399538 591690 399774
rect 591070 399454 591690 399538
rect 591070 399218 591102 399454
rect 591338 399218 591422 399454
rect 591658 399218 591690 399454
rect 591070 365774 591690 399218
rect 591070 365538 591102 365774
rect 591338 365538 591422 365774
rect 591658 365538 591690 365774
rect 591070 365454 591690 365538
rect 591070 365218 591102 365454
rect 591338 365218 591422 365454
rect 591658 365218 591690 365454
rect 591070 331774 591690 365218
rect 591070 331538 591102 331774
rect 591338 331538 591422 331774
rect 591658 331538 591690 331774
rect 591070 331454 591690 331538
rect 591070 331218 591102 331454
rect 591338 331218 591422 331454
rect 591658 331218 591690 331454
rect 591070 297774 591690 331218
rect 591070 297538 591102 297774
rect 591338 297538 591422 297774
rect 591658 297538 591690 297774
rect 591070 297454 591690 297538
rect 591070 297218 591102 297454
rect 591338 297218 591422 297454
rect 591658 297218 591690 297454
rect 591070 263774 591690 297218
rect 591070 263538 591102 263774
rect 591338 263538 591422 263774
rect 591658 263538 591690 263774
rect 591070 263454 591690 263538
rect 591070 263218 591102 263454
rect 591338 263218 591422 263454
rect 591658 263218 591690 263454
rect 591070 229774 591690 263218
rect 591070 229538 591102 229774
rect 591338 229538 591422 229774
rect 591658 229538 591690 229774
rect 591070 229454 591690 229538
rect 591070 229218 591102 229454
rect 591338 229218 591422 229454
rect 591658 229218 591690 229454
rect 591070 195774 591690 229218
rect 591070 195538 591102 195774
rect 591338 195538 591422 195774
rect 591658 195538 591690 195774
rect 591070 195454 591690 195538
rect 591070 195218 591102 195454
rect 591338 195218 591422 195454
rect 591658 195218 591690 195454
rect 591070 161774 591690 195218
rect 591070 161538 591102 161774
rect 591338 161538 591422 161774
rect 591658 161538 591690 161774
rect 591070 161454 591690 161538
rect 591070 161218 591102 161454
rect 591338 161218 591422 161454
rect 591658 161218 591690 161454
rect 591070 127774 591690 161218
rect 591070 127538 591102 127774
rect 591338 127538 591422 127774
rect 591658 127538 591690 127774
rect 591070 127454 591690 127538
rect 591070 127218 591102 127454
rect 591338 127218 591422 127454
rect 591658 127218 591690 127454
rect 591070 93774 591690 127218
rect 591070 93538 591102 93774
rect 591338 93538 591422 93774
rect 591658 93538 591690 93774
rect 591070 93454 591690 93538
rect 591070 93218 591102 93454
rect 591338 93218 591422 93454
rect 591658 93218 591690 93454
rect 591070 59774 591690 93218
rect 591070 59538 591102 59774
rect 591338 59538 591422 59774
rect 591658 59538 591690 59774
rect 591070 59454 591690 59538
rect 591070 59218 591102 59454
rect 591338 59218 591422 59454
rect 591658 59218 591690 59454
rect 591070 25774 591690 59218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 675494 592650 711002
rect 592030 675258 592062 675494
rect 592298 675258 592382 675494
rect 592618 675258 592650 675494
rect 592030 675174 592650 675258
rect 592030 674938 592062 675174
rect 592298 674938 592382 675174
rect 592618 674938 592650 675174
rect 592030 641494 592650 674938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 607494 592650 640938
rect 592030 607258 592062 607494
rect 592298 607258 592382 607494
rect 592618 607258 592650 607494
rect 592030 607174 592650 607258
rect 592030 606938 592062 607174
rect 592298 606938 592382 607174
rect 592618 606938 592650 607174
rect 592030 573494 592650 606938
rect 592030 573258 592062 573494
rect 592298 573258 592382 573494
rect 592618 573258 592650 573494
rect 592030 573174 592650 573258
rect 592030 572938 592062 573174
rect 592298 572938 592382 573174
rect 592618 572938 592650 573174
rect 592030 539494 592650 572938
rect 592030 539258 592062 539494
rect 592298 539258 592382 539494
rect 592618 539258 592650 539494
rect 592030 539174 592650 539258
rect 592030 538938 592062 539174
rect 592298 538938 592382 539174
rect 592618 538938 592650 539174
rect 592030 505494 592650 538938
rect 592030 505258 592062 505494
rect 592298 505258 592382 505494
rect 592618 505258 592650 505494
rect 592030 505174 592650 505258
rect 592030 504938 592062 505174
rect 592298 504938 592382 505174
rect 592618 504938 592650 505174
rect 592030 471494 592650 504938
rect 592030 471258 592062 471494
rect 592298 471258 592382 471494
rect 592618 471258 592650 471494
rect 592030 471174 592650 471258
rect 592030 470938 592062 471174
rect 592298 470938 592382 471174
rect 592618 470938 592650 471174
rect 592030 437494 592650 470938
rect 592030 437258 592062 437494
rect 592298 437258 592382 437494
rect 592618 437258 592650 437494
rect 592030 437174 592650 437258
rect 592030 436938 592062 437174
rect 592298 436938 592382 437174
rect 592618 436938 592650 437174
rect 592030 403494 592650 436938
rect 592030 403258 592062 403494
rect 592298 403258 592382 403494
rect 592618 403258 592650 403494
rect 592030 403174 592650 403258
rect 592030 402938 592062 403174
rect 592298 402938 592382 403174
rect 592618 402938 592650 403174
rect 592030 369494 592650 402938
rect 592030 369258 592062 369494
rect 592298 369258 592382 369494
rect 592618 369258 592650 369494
rect 592030 369174 592650 369258
rect 592030 368938 592062 369174
rect 592298 368938 592382 369174
rect 592618 368938 592650 369174
rect 592030 335494 592650 368938
rect 592030 335258 592062 335494
rect 592298 335258 592382 335494
rect 592618 335258 592650 335494
rect 592030 335174 592650 335258
rect 592030 334938 592062 335174
rect 592298 334938 592382 335174
rect 592618 334938 592650 335174
rect 592030 301494 592650 334938
rect 592030 301258 592062 301494
rect 592298 301258 592382 301494
rect 592618 301258 592650 301494
rect 592030 301174 592650 301258
rect 592030 300938 592062 301174
rect 592298 300938 592382 301174
rect 592618 300938 592650 301174
rect 592030 267494 592650 300938
rect 592030 267258 592062 267494
rect 592298 267258 592382 267494
rect 592618 267258 592650 267494
rect 592030 267174 592650 267258
rect 592030 266938 592062 267174
rect 592298 266938 592382 267174
rect 592618 266938 592650 267174
rect 592030 233494 592650 266938
rect 592030 233258 592062 233494
rect 592298 233258 592382 233494
rect 592618 233258 592650 233494
rect 592030 233174 592650 233258
rect 592030 232938 592062 233174
rect 592298 232938 592382 233174
rect 592618 232938 592650 233174
rect 592030 199494 592650 232938
rect 592030 199258 592062 199494
rect 592298 199258 592382 199494
rect 592618 199258 592650 199494
rect 592030 199174 592650 199258
rect 592030 198938 592062 199174
rect 592298 198938 592382 199174
rect 592618 198938 592650 199174
rect 592030 165494 592650 198938
rect 592030 165258 592062 165494
rect 592298 165258 592382 165494
rect 592618 165258 592650 165494
rect 592030 165174 592650 165258
rect 592030 164938 592062 165174
rect 592298 164938 592382 165174
rect 592618 164938 592650 165174
rect 592030 131494 592650 164938
rect 592030 131258 592062 131494
rect 592298 131258 592382 131494
rect 592618 131258 592650 131494
rect 592030 131174 592650 131258
rect 592030 130938 592062 131174
rect 592298 130938 592382 131174
rect 592618 130938 592650 131174
rect 592030 97494 592650 130938
rect 592030 97258 592062 97494
rect 592298 97258 592382 97494
rect 592618 97258 592650 97494
rect 592030 97174 592650 97258
rect 592030 96938 592062 97174
rect 592298 96938 592382 97174
rect 592618 96938 592650 97174
rect 592030 63494 592650 96938
rect 592030 63258 592062 63494
rect 592298 63258 592382 63494
rect 592618 63258 592650 63494
rect 592030 63174 592650 63258
rect 592030 62938 592062 63174
rect 592298 62938 592382 63174
rect 592618 62938 592650 63174
rect 592030 29494 592650 62938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 675258 -8458 675494
rect -8374 675258 -8138 675494
rect -8694 674938 -8458 675174
rect -8374 674938 -8138 675174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 607258 -8458 607494
rect -8374 607258 -8138 607494
rect -8694 606938 -8458 607174
rect -8374 606938 -8138 607174
rect -8694 573258 -8458 573494
rect -8374 573258 -8138 573494
rect -8694 572938 -8458 573174
rect -8374 572938 -8138 573174
rect -8694 539258 -8458 539494
rect -8374 539258 -8138 539494
rect -8694 538938 -8458 539174
rect -8374 538938 -8138 539174
rect -8694 505258 -8458 505494
rect -8374 505258 -8138 505494
rect -8694 504938 -8458 505174
rect -8374 504938 -8138 505174
rect -8694 471258 -8458 471494
rect -8374 471258 -8138 471494
rect -8694 470938 -8458 471174
rect -8374 470938 -8138 471174
rect -8694 437258 -8458 437494
rect -8374 437258 -8138 437494
rect -8694 436938 -8458 437174
rect -8374 436938 -8138 437174
rect -8694 403258 -8458 403494
rect -8374 403258 -8138 403494
rect -8694 402938 -8458 403174
rect -8374 402938 -8138 403174
rect -8694 369258 -8458 369494
rect -8374 369258 -8138 369494
rect -8694 368938 -8458 369174
rect -8374 368938 -8138 369174
rect -8694 335258 -8458 335494
rect -8374 335258 -8138 335494
rect -8694 334938 -8458 335174
rect -8374 334938 -8138 335174
rect -8694 301258 -8458 301494
rect -8374 301258 -8138 301494
rect -8694 300938 -8458 301174
rect -8374 300938 -8138 301174
rect -8694 267258 -8458 267494
rect -8374 267258 -8138 267494
rect -8694 266938 -8458 267174
rect -8374 266938 -8138 267174
rect -8694 233258 -8458 233494
rect -8374 233258 -8138 233494
rect -8694 232938 -8458 233174
rect -8374 232938 -8138 233174
rect -8694 199258 -8458 199494
rect -8374 199258 -8138 199494
rect -8694 198938 -8458 199174
rect -8374 198938 -8138 199174
rect -8694 165258 -8458 165494
rect -8374 165258 -8138 165494
rect -8694 164938 -8458 165174
rect -8374 164938 -8138 165174
rect -8694 131258 -8458 131494
rect -8374 131258 -8138 131494
rect -8694 130938 -8458 131174
rect -8374 130938 -8138 131174
rect -8694 97258 -8458 97494
rect -8374 97258 -8138 97494
rect -8694 96938 -8458 97174
rect -8374 96938 -8138 97174
rect -8694 63258 -8458 63494
rect -8374 63258 -8138 63494
rect -8694 62938 -8458 63174
rect -8374 62938 -8138 63174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 671538 -7498 671774
rect -7414 671538 -7178 671774
rect -7734 671218 -7498 671454
rect -7414 671218 -7178 671454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 603538 -7498 603774
rect -7414 603538 -7178 603774
rect -7734 603218 -7498 603454
rect -7414 603218 -7178 603454
rect -7734 569538 -7498 569774
rect -7414 569538 -7178 569774
rect -7734 569218 -7498 569454
rect -7414 569218 -7178 569454
rect -7734 535538 -7498 535774
rect -7414 535538 -7178 535774
rect -7734 535218 -7498 535454
rect -7414 535218 -7178 535454
rect -7734 501538 -7498 501774
rect -7414 501538 -7178 501774
rect -7734 501218 -7498 501454
rect -7414 501218 -7178 501454
rect -7734 467538 -7498 467774
rect -7414 467538 -7178 467774
rect -7734 467218 -7498 467454
rect -7414 467218 -7178 467454
rect -7734 433538 -7498 433774
rect -7414 433538 -7178 433774
rect -7734 433218 -7498 433454
rect -7414 433218 -7178 433454
rect -7734 399538 -7498 399774
rect -7414 399538 -7178 399774
rect -7734 399218 -7498 399454
rect -7414 399218 -7178 399454
rect -7734 365538 -7498 365774
rect -7414 365538 -7178 365774
rect -7734 365218 -7498 365454
rect -7414 365218 -7178 365454
rect -7734 331538 -7498 331774
rect -7414 331538 -7178 331774
rect -7734 331218 -7498 331454
rect -7414 331218 -7178 331454
rect -7734 297538 -7498 297774
rect -7414 297538 -7178 297774
rect -7734 297218 -7498 297454
rect -7414 297218 -7178 297454
rect -7734 263538 -7498 263774
rect -7414 263538 -7178 263774
rect -7734 263218 -7498 263454
rect -7414 263218 -7178 263454
rect -7734 229538 -7498 229774
rect -7414 229538 -7178 229774
rect -7734 229218 -7498 229454
rect -7414 229218 -7178 229454
rect -7734 195538 -7498 195774
rect -7414 195538 -7178 195774
rect -7734 195218 -7498 195454
rect -7414 195218 -7178 195454
rect -7734 161538 -7498 161774
rect -7414 161538 -7178 161774
rect -7734 161218 -7498 161454
rect -7414 161218 -7178 161454
rect -7734 127538 -7498 127774
rect -7414 127538 -7178 127774
rect -7734 127218 -7498 127454
rect -7414 127218 -7178 127454
rect -7734 93538 -7498 93774
rect -7414 93538 -7178 93774
rect -7734 93218 -7498 93454
rect -7414 93218 -7178 93454
rect -7734 59538 -7498 59774
rect -7414 59538 -7178 59774
rect -7734 59218 -7498 59454
rect -7414 59218 -7178 59454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 667818 -6538 668054
rect -6454 667818 -6218 668054
rect -6774 667498 -6538 667734
rect -6454 667498 -6218 667734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 599818 -6538 600054
rect -6454 599818 -6218 600054
rect -6774 599498 -6538 599734
rect -6454 599498 -6218 599734
rect -6774 565818 -6538 566054
rect -6454 565818 -6218 566054
rect -6774 565498 -6538 565734
rect -6454 565498 -6218 565734
rect -6774 531818 -6538 532054
rect -6454 531818 -6218 532054
rect -6774 531498 -6538 531734
rect -6454 531498 -6218 531734
rect -6774 497818 -6538 498054
rect -6454 497818 -6218 498054
rect -6774 497498 -6538 497734
rect -6454 497498 -6218 497734
rect -6774 463818 -6538 464054
rect -6454 463818 -6218 464054
rect -6774 463498 -6538 463734
rect -6454 463498 -6218 463734
rect -6774 429818 -6538 430054
rect -6454 429818 -6218 430054
rect -6774 429498 -6538 429734
rect -6454 429498 -6218 429734
rect -6774 395818 -6538 396054
rect -6454 395818 -6218 396054
rect -6774 395498 -6538 395734
rect -6454 395498 -6218 395734
rect -6774 361818 -6538 362054
rect -6454 361818 -6218 362054
rect -6774 361498 -6538 361734
rect -6454 361498 -6218 361734
rect -6774 327818 -6538 328054
rect -6454 327818 -6218 328054
rect -6774 327498 -6538 327734
rect -6454 327498 -6218 327734
rect -6774 293818 -6538 294054
rect -6454 293818 -6218 294054
rect -6774 293498 -6538 293734
rect -6454 293498 -6218 293734
rect -6774 259818 -6538 260054
rect -6454 259818 -6218 260054
rect -6774 259498 -6538 259734
rect -6454 259498 -6218 259734
rect -6774 225818 -6538 226054
rect -6454 225818 -6218 226054
rect -6774 225498 -6538 225734
rect -6454 225498 -6218 225734
rect -6774 191818 -6538 192054
rect -6454 191818 -6218 192054
rect -6774 191498 -6538 191734
rect -6454 191498 -6218 191734
rect -6774 157818 -6538 158054
rect -6454 157818 -6218 158054
rect -6774 157498 -6538 157734
rect -6454 157498 -6218 157734
rect -6774 123818 -6538 124054
rect -6454 123818 -6218 124054
rect -6774 123498 -6538 123734
rect -6454 123498 -6218 123734
rect -6774 89818 -6538 90054
rect -6454 89818 -6218 90054
rect -6774 89498 -6538 89734
rect -6454 89498 -6218 89734
rect -6774 55818 -6538 56054
rect -6454 55818 -6218 56054
rect -6774 55498 -6538 55734
rect -6454 55498 -6218 55734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 698098 -5578 698334
rect -5494 698098 -5258 698334
rect -5814 697778 -5578 698014
rect -5494 697778 -5258 698014
rect -5814 664098 -5578 664334
rect -5494 664098 -5258 664334
rect -5814 663778 -5578 664014
rect -5494 663778 -5258 664014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 596098 -5578 596334
rect -5494 596098 -5258 596334
rect -5814 595778 -5578 596014
rect -5494 595778 -5258 596014
rect -5814 562098 -5578 562334
rect -5494 562098 -5258 562334
rect -5814 561778 -5578 562014
rect -5494 561778 -5258 562014
rect -5814 528098 -5578 528334
rect -5494 528098 -5258 528334
rect -5814 527778 -5578 528014
rect -5494 527778 -5258 528014
rect -5814 494098 -5578 494334
rect -5494 494098 -5258 494334
rect -5814 493778 -5578 494014
rect -5494 493778 -5258 494014
rect -5814 460098 -5578 460334
rect -5494 460098 -5258 460334
rect -5814 459778 -5578 460014
rect -5494 459778 -5258 460014
rect -5814 426098 -5578 426334
rect -5494 426098 -5258 426334
rect -5814 425778 -5578 426014
rect -5494 425778 -5258 426014
rect -5814 392098 -5578 392334
rect -5494 392098 -5258 392334
rect -5814 391778 -5578 392014
rect -5494 391778 -5258 392014
rect -5814 358098 -5578 358334
rect -5494 358098 -5258 358334
rect -5814 357778 -5578 358014
rect -5494 357778 -5258 358014
rect -5814 324098 -5578 324334
rect -5494 324098 -5258 324334
rect -5814 323778 -5578 324014
rect -5494 323778 -5258 324014
rect -5814 290098 -5578 290334
rect -5494 290098 -5258 290334
rect -5814 289778 -5578 290014
rect -5494 289778 -5258 290014
rect -5814 256098 -5578 256334
rect -5494 256098 -5258 256334
rect -5814 255778 -5578 256014
rect -5494 255778 -5258 256014
rect -5814 222098 -5578 222334
rect -5494 222098 -5258 222334
rect -5814 221778 -5578 222014
rect -5494 221778 -5258 222014
rect -5814 188098 -5578 188334
rect -5494 188098 -5258 188334
rect -5814 187778 -5578 188014
rect -5494 187778 -5258 188014
rect -5814 154098 -5578 154334
rect -5494 154098 -5258 154334
rect -5814 153778 -5578 154014
rect -5494 153778 -5258 154014
rect -5814 120098 -5578 120334
rect -5494 120098 -5258 120334
rect -5814 119778 -5578 120014
rect -5494 119778 -5258 120014
rect -5814 86098 -5578 86334
rect -5494 86098 -5258 86334
rect -5814 85778 -5578 86014
rect -5494 85778 -5258 86014
rect -5814 52098 -5578 52334
rect -5494 52098 -5258 52334
rect -5814 51778 -5578 52014
rect -5494 51778 -5258 52014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 694378 -4618 694614
rect -4534 694378 -4298 694614
rect -4854 694058 -4618 694294
rect -4534 694058 -4298 694294
rect -4854 660378 -4618 660614
rect -4534 660378 -4298 660614
rect -4854 660058 -4618 660294
rect -4534 660058 -4298 660294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 592378 -4618 592614
rect -4534 592378 -4298 592614
rect -4854 592058 -4618 592294
rect -4534 592058 -4298 592294
rect -4854 558378 -4618 558614
rect -4534 558378 -4298 558614
rect -4854 558058 -4618 558294
rect -4534 558058 -4298 558294
rect -4854 524378 -4618 524614
rect -4534 524378 -4298 524614
rect -4854 524058 -4618 524294
rect -4534 524058 -4298 524294
rect -4854 490378 -4618 490614
rect -4534 490378 -4298 490614
rect -4854 490058 -4618 490294
rect -4534 490058 -4298 490294
rect -4854 456378 -4618 456614
rect -4534 456378 -4298 456614
rect -4854 456058 -4618 456294
rect -4534 456058 -4298 456294
rect -4854 422378 -4618 422614
rect -4534 422378 -4298 422614
rect -4854 422058 -4618 422294
rect -4534 422058 -4298 422294
rect -4854 388378 -4618 388614
rect -4534 388378 -4298 388614
rect -4854 388058 -4618 388294
rect -4534 388058 -4298 388294
rect -4854 354378 -4618 354614
rect -4534 354378 -4298 354614
rect -4854 354058 -4618 354294
rect -4534 354058 -4298 354294
rect -4854 320378 -4618 320614
rect -4534 320378 -4298 320614
rect -4854 320058 -4618 320294
rect -4534 320058 -4298 320294
rect -4854 286378 -4618 286614
rect -4534 286378 -4298 286614
rect -4854 286058 -4618 286294
rect -4534 286058 -4298 286294
rect -4854 252378 -4618 252614
rect -4534 252378 -4298 252614
rect -4854 252058 -4618 252294
rect -4534 252058 -4298 252294
rect -4854 218378 -4618 218614
rect -4534 218378 -4298 218614
rect -4854 218058 -4618 218294
rect -4534 218058 -4298 218294
rect -4854 184378 -4618 184614
rect -4534 184378 -4298 184614
rect -4854 184058 -4618 184294
rect -4534 184058 -4298 184294
rect -4854 150378 -4618 150614
rect -4534 150378 -4298 150614
rect -4854 150058 -4618 150294
rect -4534 150058 -4298 150294
rect -4854 116378 -4618 116614
rect -4534 116378 -4298 116614
rect -4854 116058 -4618 116294
rect -4534 116058 -4298 116294
rect -4854 82378 -4618 82614
rect -4534 82378 -4298 82614
rect -4854 82058 -4618 82294
rect -4534 82058 -4298 82294
rect -4854 48378 -4618 48614
rect -4534 48378 -4298 48614
rect -4854 48058 -4618 48294
rect -4534 48058 -4298 48294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 690658 -3658 690894
rect -3574 690658 -3338 690894
rect -3894 690338 -3658 690574
rect -3574 690338 -3338 690574
rect -3894 656658 -3658 656894
rect -3574 656658 -3338 656894
rect -3894 656338 -3658 656574
rect -3574 656338 -3338 656574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 588658 -3658 588894
rect -3574 588658 -3338 588894
rect -3894 588338 -3658 588574
rect -3574 588338 -3338 588574
rect -3894 554658 -3658 554894
rect -3574 554658 -3338 554894
rect -3894 554338 -3658 554574
rect -3574 554338 -3338 554574
rect -3894 520658 -3658 520894
rect -3574 520658 -3338 520894
rect -3894 520338 -3658 520574
rect -3574 520338 -3338 520574
rect -3894 486658 -3658 486894
rect -3574 486658 -3338 486894
rect -3894 486338 -3658 486574
rect -3574 486338 -3338 486574
rect -3894 452658 -3658 452894
rect -3574 452658 -3338 452894
rect -3894 452338 -3658 452574
rect -3574 452338 -3338 452574
rect -3894 418658 -3658 418894
rect -3574 418658 -3338 418894
rect -3894 418338 -3658 418574
rect -3574 418338 -3338 418574
rect -3894 384658 -3658 384894
rect -3574 384658 -3338 384894
rect -3894 384338 -3658 384574
rect -3574 384338 -3338 384574
rect -3894 350658 -3658 350894
rect -3574 350658 -3338 350894
rect -3894 350338 -3658 350574
rect -3574 350338 -3338 350574
rect -3894 316658 -3658 316894
rect -3574 316658 -3338 316894
rect -3894 316338 -3658 316574
rect -3574 316338 -3338 316574
rect -3894 282658 -3658 282894
rect -3574 282658 -3338 282894
rect -3894 282338 -3658 282574
rect -3574 282338 -3338 282574
rect -3894 248658 -3658 248894
rect -3574 248658 -3338 248894
rect -3894 248338 -3658 248574
rect -3574 248338 -3338 248574
rect -3894 214658 -3658 214894
rect -3574 214658 -3338 214894
rect -3894 214338 -3658 214574
rect -3574 214338 -3338 214574
rect -3894 180658 -3658 180894
rect -3574 180658 -3338 180894
rect -3894 180338 -3658 180574
rect -3574 180338 -3338 180574
rect -3894 146658 -3658 146894
rect -3574 146658 -3338 146894
rect -3894 146338 -3658 146574
rect -3574 146338 -3338 146574
rect -3894 112658 -3658 112894
rect -3574 112658 -3338 112894
rect -3894 112338 -3658 112574
rect -3574 112338 -3338 112574
rect -3894 78658 -3658 78894
rect -3574 78658 -3338 78894
rect -3894 78338 -3658 78574
rect -3574 78338 -3338 78574
rect -3894 44658 -3658 44894
rect -3574 44658 -3338 44894
rect -3894 44338 -3658 44574
rect -3574 44338 -3338 44574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 686938 -2698 687174
rect -2614 686938 -2378 687174
rect -2934 686618 -2698 686854
rect -2614 686618 -2378 686854
rect -2934 652938 -2698 653174
rect -2614 652938 -2378 653174
rect -2934 652618 -2698 652854
rect -2614 652618 -2378 652854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 584938 -2698 585174
rect -2614 584938 -2378 585174
rect -2934 584618 -2698 584854
rect -2614 584618 -2378 584854
rect -2934 550938 -2698 551174
rect -2614 550938 -2378 551174
rect -2934 550618 -2698 550854
rect -2614 550618 -2378 550854
rect -2934 516938 -2698 517174
rect -2614 516938 -2378 517174
rect -2934 516618 -2698 516854
rect -2614 516618 -2378 516854
rect -2934 482938 -2698 483174
rect -2614 482938 -2378 483174
rect -2934 482618 -2698 482854
rect -2614 482618 -2378 482854
rect -2934 448938 -2698 449174
rect -2614 448938 -2378 449174
rect -2934 448618 -2698 448854
rect -2614 448618 -2378 448854
rect -2934 414938 -2698 415174
rect -2614 414938 -2378 415174
rect -2934 414618 -2698 414854
rect -2614 414618 -2378 414854
rect -2934 380938 -2698 381174
rect -2614 380938 -2378 381174
rect -2934 380618 -2698 380854
rect -2614 380618 -2378 380854
rect -2934 346938 -2698 347174
rect -2614 346938 -2378 347174
rect -2934 346618 -2698 346854
rect -2614 346618 -2378 346854
rect -2934 312938 -2698 313174
rect -2614 312938 -2378 313174
rect -2934 312618 -2698 312854
rect -2614 312618 -2378 312854
rect -2934 278938 -2698 279174
rect -2614 278938 -2378 279174
rect -2934 278618 -2698 278854
rect -2614 278618 -2378 278854
rect -2934 244938 -2698 245174
rect -2614 244938 -2378 245174
rect -2934 244618 -2698 244854
rect -2614 244618 -2378 244854
rect -2934 210938 -2698 211174
rect -2614 210938 -2378 211174
rect -2934 210618 -2698 210854
rect -2614 210618 -2378 210854
rect -2934 176938 -2698 177174
rect -2614 176938 -2378 177174
rect -2934 176618 -2698 176854
rect -2614 176618 -2378 176854
rect -2934 142938 -2698 143174
rect -2614 142938 -2378 143174
rect -2934 142618 -2698 142854
rect -2614 142618 -2378 142854
rect -2934 108938 -2698 109174
rect -2614 108938 -2378 109174
rect -2934 108618 -2698 108854
rect -2614 108618 -2378 108854
rect -2934 74938 -2698 75174
rect -2614 74938 -2378 75174
rect -2934 74618 -2698 74854
rect -2614 74618 -2378 74854
rect -2934 40938 -2698 41174
rect -2614 40938 -2378 41174
rect -2934 40618 -2698 40854
rect -2614 40618 -2378 40854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 683218 -1738 683454
rect -1654 683218 -1418 683454
rect -1974 682898 -1738 683134
rect -1654 682898 -1418 683134
rect -1974 649218 -1738 649454
rect -1654 649218 -1418 649454
rect -1974 648898 -1738 649134
rect -1654 648898 -1418 649134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 581218 -1738 581454
rect -1654 581218 -1418 581454
rect -1974 580898 -1738 581134
rect -1654 580898 -1418 581134
rect -1974 547218 -1738 547454
rect -1654 547218 -1418 547454
rect -1974 546898 -1738 547134
rect -1654 546898 -1418 547134
rect -1974 513218 -1738 513454
rect -1654 513218 -1418 513454
rect -1974 512898 -1738 513134
rect -1654 512898 -1418 513134
rect -1974 479218 -1738 479454
rect -1654 479218 -1418 479454
rect -1974 478898 -1738 479134
rect -1654 478898 -1418 479134
rect -1974 445218 -1738 445454
rect -1654 445218 -1418 445454
rect -1974 444898 -1738 445134
rect -1654 444898 -1418 445134
rect -1974 411218 -1738 411454
rect -1654 411218 -1418 411454
rect -1974 410898 -1738 411134
rect -1654 410898 -1418 411134
rect -1974 377218 -1738 377454
rect -1654 377218 -1418 377454
rect -1974 376898 -1738 377134
rect -1654 376898 -1418 377134
rect -1974 343218 -1738 343454
rect -1654 343218 -1418 343454
rect -1974 342898 -1738 343134
rect -1654 342898 -1418 343134
rect -1974 309218 -1738 309454
rect -1654 309218 -1418 309454
rect -1974 308898 -1738 309134
rect -1654 308898 -1418 309134
rect -1974 275218 -1738 275454
rect -1654 275218 -1418 275454
rect -1974 274898 -1738 275134
rect -1654 274898 -1418 275134
rect -1974 241218 -1738 241454
rect -1654 241218 -1418 241454
rect -1974 240898 -1738 241134
rect -1654 240898 -1418 241134
rect -1974 207218 -1738 207454
rect -1654 207218 -1418 207454
rect -1974 206898 -1738 207134
rect -1654 206898 -1418 207134
rect -1974 173218 -1738 173454
rect -1654 173218 -1418 173454
rect -1974 172898 -1738 173134
rect -1654 172898 -1418 173134
rect -1974 139218 -1738 139454
rect -1654 139218 -1418 139454
rect -1974 138898 -1738 139134
rect -1654 138898 -1418 139134
rect -1974 105218 -1738 105454
rect -1654 105218 -1418 105454
rect -1974 104898 -1738 105134
rect -1654 104898 -1418 105134
rect -1974 71218 -1738 71454
rect -1654 71218 -1418 71454
rect -1974 70898 -1738 71134
rect -1654 70898 -1418 71134
rect -1974 37218 -1738 37454
rect -1654 37218 -1418 37454
rect -1974 36898 -1738 37134
rect -1654 36898 -1418 37134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 683218 2062 683454
rect 2146 683218 2382 683454
rect 1826 682898 2062 683134
rect 2146 682898 2382 683134
rect 1826 649218 2062 649454
rect 2146 649218 2382 649454
rect 1826 648898 2062 649134
rect 2146 648898 2382 649134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 581218 2062 581454
rect 2146 581218 2382 581454
rect 1826 580898 2062 581134
rect 2146 580898 2382 581134
rect 1826 547218 2062 547454
rect 2146 547218 2382 547454
rect 1826 546898 2062 547134
rect 2146 546898 2382 547134
rect 1826 513218 2062 513454
rect 2146 513218 2382 513454
rect 1826 512898 2062 513134
rect 2146 512898 2382 513134
rect 1826 479218 2062 479454
rect 2146 479218 2382 479454
rect 1826 478898 2062 479134
rect 2146 478898 2382 479134
rect 1826 445218 2062 445454
rect 2146 445218 2382 445454
rect 1826 444898 2062 445134
rect 2146 444898 2382 445134
rect 1826 411218 2062 411454
rect 2146 411218 2382 411454
rect 1826 410898 2062 411134
rect 2146 410898 2382 411134
rect 1826 377218 2062 377454
rect 2146 377218 2382 377454
rect 1826 376898 2062 377134
rect 2146 376898 2382 377134
rect 1826 343218 2062 343454
rect 2146 343218 2382 343454
rect 1826 342898 2062 343134
rect 2146 342898 2382 343134
rect 1826 309218 2062 309454
rect 2146 309218 2382 309454
rect 1826 308898 2062 309134
rect 2146 308898 2382 309134
rect 1826 275218 2062 275454
rect 2146 275218 2382 275454
rect 1826 274898 2062 275134
rect 2146 274898 2382 275134
rect 1826 241218 2062 241454
rect 2146 241218 2382 241454
rect 1826 240898 2062 241134
rect 2146 240898 2382 241134
rect 1826 207218 2062 207454
rect 2146 207218 2382 207454
rect 1826 206898 2062 207134
rect 2146 206898 2382 207134
rect 1826 173218 2062 173454
rect 2146 173218 2382 173454
rect 1826 172898 2062 173134
rect 2146 172898 2382 173134
rect 1826 139218 2062 139454
rect 2146 139218 2382 139454
rect 1826 138898 2062 139134
rect 2146 138898 2382 139134
rect 1826 105218 2062 105454
rect 2146 105218 2382 105454
rect 1826 104898 2062 105134
rect 2146 104898 2382 105134
rect 1826 71218 2062 71454
rect 2146 71218 2382 71454
rect 1826 70898 2062 71134
rect 2146 70898 2382 71134
rect 1826 37218 2062 37454
rect 2146 37218 2382 37454
rect 1826 36898 2062 37134
rect 2146 36898 2382 37134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 686938 5782 687174
rect 5866 686938 6102 687174
rect 5546 686618 5782 686854
rect 5866 686618 6102 686854
rect 5546 652938 5782 653174
rect 5866 652938 6102 653174
rect 5546 652618 5782 652854
rect 5866 652618 6102 652854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 584938 5782 585174
rect 5866 584938 6102 585174
rect 5546 584618 5782 584854
rect 5866 584618 6102 584854
rect 5546 550938 5782 551174
rect 5866 550938 6102 551174
rect 5546 550618 5782 550854
rect 5866 550618 6102 550854
rect 5546 516938 5782 517174
rect 5866 516938 6102 517174
rect 5546 516618 5782 516854
rect 5866 516618 6102 516854
rect 5546 482938 5782 483174
rect 5866 482938 6102 483174
rect 5546 482618 5782 482854
rect 5866 482618 6102 482854
rect 5546 448938 5782 449174
rect 5866 448938 6102 449174
rect 5546 448618 5782 448854
rect 5866 448618 6102 448854
rect 5546 414938 5782 415174
rect 5866 414938 6102 415174
rect 5546 414618 5782 414854
rect 5866 414618 6102 414854
rect 5546 380938 5782 381174
rect 5866 380938 6102 381174
rect 5546 380618 5782 380854
rect 5866 380618 6102 380854
rect 5546 346938 5782 347174
rect 5866 346938 6102 347174
rect 5546 346618 5782 346854
rect 5866 346618 6102 346854
rect 5546 312938 5782 313174
rect 5866 312938 6102 313174
rect 5546 312618 5782 312854
rect 5866 312618 6102 312854
rect 5546 278938 5782 279174
rect 5866 278938 6102 279174
rect 5546 278618 5782 278854
rect 5866 278618 6102 278854
rect 5546 244938 5782 245174
rect 5866 244938 6102 245174
rect 5546 244618 5782 244854
rect 5866 244618 6102 244854
rect 5546 210938 5782 211174
rect 5866 210938 6102 211174
rect 5546 210618 5782 210854
rect 5866 210618 6102 210854
rect 5546 176938 5782 177174
rect 5866 176938 6102 177174
rect 5546 176618 5782 176854
rect 5866 176618 6102 176854
rect 5546 142938 5782 143174
rect 5866 142938 6102 143174
rect 5546 142618 5782 142854
rect 5866 142618 6102 142854
rect 5546 108938 5782 109174
rect 5866 108938 6102 109174
rect 5546 108618 5782 108854
rect 5866 108618 6102 108854
rect 5546 74938 5782 75174
rect 5866 74938 6102 75174
rect 5546 74618 5782 74854
rect 5866 74618 6102 74854
rect 5546 40938 5782 41174
rect 5866 40938 6102 41174
rect 5546 40618 5782 40854
rect 5866 40618 6102 40854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 690658 9502 690894
rect 9586 690658 9822 690894
rect 9266 690338 9502 690574
rect 9586 690338 9822 690574
rect 9266 656658 9502 656894
rect 9586 656658 9822 656894
rect 9266 656338 9502 656574
rect 9586 656338 9822 656574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 588658 9502 588894
rect 9586 588658 9822 588894
rect 9266 588338 9502 588574
rect 9586 588338 9822 588574
rect 9266 554658 9502 554894
rect 9586 554658 9822 554894
rect 9266 554338 9502 554574
rect 9586 554338 9822 554574
rect 9266 520658 9502 520894
rect 9586 520658 9822 520894
rect 9266 520338 9502 520574
rect 9586 520338 9822 520574
rect 9266 486658 9502 486894
rect 9586 486658 9822 486894
rect 9266 486338 9502 486574
rect 9586 486338 9822 486574
rect 9266 452658 9502 452894
rect 9586 452658 9822 452894
rect 9266 452338 9502 452574
rect 9586 452338 9822 452574
rect 9266 418658 9502 418894
rect 9586 418658 9822 418894
rect 9266 418338 9502 418574
rect 9586 418338 9822 418574
rect 9266 384658 9502 384894
rect 9586 384658 9822 384894
rect 9266 384338 9502 384574
rect 9586 384338 9822 384574
rect 9266 350658 9502 350894
rect 9586 350658 9822 350894
rect 9266 350338 9502 350574
rect 9586 350338 9822 350574
rect 9266 316658 9502 316894
rect 9586 316658 9822 316894
rect 9266 316338 9502 316574
rect 9586 316338 9822 316574
rect 9266 282658 9502 282894
rect 9586 282658 9822 282894
rect 9266 282338 9502 282574
rect 9586 282338 9822 282574
rect 9266 248658 9502 248894
rect 9586 248658 9822 248894
rect 9266 248338 9502 248574
rect 9586 248338 9822 248574
rect 9266 214658 9502 214894
rect 9586 214658 9822 214894
rect 9266 214338 9502 214574
rect 9586 214338 9822 214574
rect 9266 180658 9502 180894
rect 9586 180658 9822 180894
rect 9266 180338 9502 180574
rect 9586 180338 9822 180574
rect 9266 146658 9502 146894
rect 9586 146658 9822 146894
rect 9266 146338 9502 146574
rect 9586 146338 9822 146574
rect 9266 112658 9502 112894
rect 9586 112658 9822 112894
rect 9266 112338 9502 112574
rect 9586 112338 9822 112574
rect 9266 78658 9502 78894
rect 9586 78658 9822 78894
rect 9266 78338 9502 78574
rect 9586 78338 9822 78574
rect 9266 44658 9502 44894
rect 9586 44658 9822 44894
rect 9266 44338 9502 44574
rect 9586 44338 9822 44574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 694378 13222 694614
rect 13306 694378 13542 694614
rect 12986 694058 13222 694294
rect 13306 694058 13542 694294
rect 12986 660378 13222 660614
rect 13306 660378 13542 660614
rect 12986 660058 13222 660294
rect 13306 660058 13542 660294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 592378 13222 592614
rect 13306 592378 13542 592614
rect 12986 592058 13222 592294
rect 13306 592058 13542 592294
rect 12986 558378 13222 558614
rect 13306 558378 13542 558614
rect 12986 558058 13222 558294
rect 13306 558058 13542 558294
rect 12986 524378 13222 524614
rect 13306 524378 13542 524614
rect 12986 524058 13222 524294
rect 13306 524058 13542 524294
rect 12986 490378 13222 490614
rect 13306 490378 13542 490614
rect 12986 490058 13222 490294
rect 13306 490058 13542 490294
rect 12986 456378 13222 456614
rect 13306 456378 13542 456614
rect 12986 456058 13222 456294
rect 13306 456058 13542 456294
rect 12986 422378 13222 422614
rect 13306 422378 13542 422614
rect 12986 422058 13222 422294
rect 13306 422058 13542 422294
rect 12986 388378 13222 388614
rect 13306 388378 13542 388614
rect 12986 388058 13222 388294
rect 13306 388058 13542 388294
rect 12986 354378 13222 354614
rect 13306 354378 13542 354614
rect 12986 354058 13222 354294
rect 13306 354058 13542 354294
rect 12986 320378 13222 320614
rect 13306 320378 13542 320614
rect 12986 320058 13222 320294
rect 13306 320058 13542 320294
rect 12986 286378 13222 286614
rect 13306 286378 13542 286614
rect 12986 286058 13222 286294
rect 13306 286058 13542 286294
rect 12986 252378 13222 252614
rect 13306 252378 13542 252614
rect 12986 252058 13222 252294
rect 13306 252058 13542 252294
rect 12986 218378 13222 218614
rect 13306 218378 13542 218614
rect 12986 218058 13222 218294
rect 13306 218058 13542 218294
rect 12986 184378 13222 184614
rect 13306 184378 13542 184614
rect 12986 184058 13222 184294
rect 13306 184058 13542 184294
rect 12986 150378 13222 150614
rect 13306 150378 13542 150614
rect 12986 150058 13222 150294
rect 13306 150058 13542 150294
rect 12986 116378 13222 116614
rect 13306 116378 13542 116614
rect 12986 116058 13222 116294
rect 13306 116058 13542 116294
rect 12986 82378 13222 82614
rect 13306 82378 13542 82614
rect 12986 82058 13222 82294
rect 13306 82058 13542 82294
rect 12986 48378 13222 48614
rect 13306 48378 13542 48614
rect 12986 48058 13222 48294
rect 13306 48058 13542 48294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 698098 16942 698334
rect 17026 698098 17262 698334
rect 16706 697778 16942 698014
rect 17026 697778 17262 698014
rect 16706 664098 16942 664334
rect 17026 664098 17262 664334
rect 16706 663778 16942 664014
rect 17026 663778 17262 664014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 596098 16942 596334
rect 17026 596098 17262 596334
rect 16706 595778 16942 596014
rect 17026 595778 17262 596014
rect 16706 562098 16942 562334
rect 17026 562098 17262 562334
rect 16706 561778 16942 562014
rect 17026 561778 17262 562014
rect 16706 528098 16942 528334
rect 17026 528098 17262 528334
rect 16706 527778 16942 528014
rect 17026 527778 17262 528014
rect 16706 494098 16942 494334
rect 17026 494098 17262 494334
rect 16706 493778 16942 494014
rect 17026 493778 17262 494014
rect 16706 460098 16942 460334
rect 17026 460098 17262 460334
rect 16706 459778 16942 460014
rect 17026 459778 17262 460014
rect 16706 426098 16942 426334
rect 17026 426098 17262 426334
rect 16706 425778 16942 426014
rect 17026 425778 17262 426014
rect 16706 392098 16942 392334
rect 17026 392098 17262 392334
rect 16706 391778 16942 392014
rect 17026 391778 17262 392014
rect 16706 358098 16942 358334
rect 17026 358098 17262 358334
rect 16706 357778 16942 358014
rect 17026 357778 17262 358014
rect 16706 324098 16942 324334
rect 17026 324098 17262 324334
rect 16706 323778 16942 324014
rect 17026 323778 17262 324014
rect 16706 290098 16942 290334
rect 17026 290098 17262 290334
rect 16706 289778 16942 290014
rect 17026 289778 17262 290014
rect 16706 256098 16942 256334
rect 17026 256098 17262 256334
rect 16706 255778 16942 256014
rect 17026 255778 17262 256014
rect 16706 222098 16942 222334
rect 17026 222098 17262 222334
rect 16706 221778 16942 222014
rect 17026 221778 17262 222014
rect 16706 188098 16942 188334
rect 17026 188098 17262 188334
rect 16706 187778 16942 188014
rect 17026 187778 17262 188014
rect 16706 154098 16942 154334
rect 17026 154098 17262 154334
rect 16706 153778 16942 154014
rect 17026 153778 17262 154014
rect 16706 120098 16942 120334
rect 17026 120098 17262 120334
rect 16706 119778 16942 120014
rect 17026 119778 17262 120014
rect 16706 86098 16942 86334
rect 17026 86098 17262 86334
rect 16706 85778 16942 86014
rect 17026 85778 17262 86014
rect 16706 52098 16942 52334
rect 17026 52098 17262 52334
rect 16706 51778 16942 52014
rect 17026 51778 17262 52014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 667818 20662 668054
rect 20746 667818 20982 668054
rect 20426 667498 20662 667734
rect 20746 667498 20982 667734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 599818 20662 600054
rect 20746 599818 20982 600054
rect 20426 599498 20662 599734
rect 20746 599498 20982 599734
rect 20426 565818 20662 566054
rect 20746 565818 20982 566054
rect 20426 565498 20662 565734
rect 20746 565498 20982 565734
rect 20426 531818 20662 532054
rect 20746 531818 20982 532054
rect 20426 531498 20662 531734
rect 20746 531498 20982 531734
rect 20426 497818 20662 498054
rect 20746 497818 20982 498054
rect 20426 497498 20662 497734
rect 20746 497498 20982 497734
rect 20426 463818 20662 464054
rect 20746 463818 20982 464054
rect 20426 463498 20662 463734
rect 20746 463498 20982 463734
rect 20426 429818 20662 430054
rect 20746 429818 20982 430054
rect 20426 429498 20662 429734
rect 20746 429498 20982 429734
rect 20426 395818 20662 396054
rect 20746 395818 20982 396054
rect 20426 395498 20662 395734
rect 20746 395498 20982 395734
rect 20426 361818 20662 362054
rect 20746 361818 20982 362054
rect 20426 361498 20662 361734
rect 20746 361498 20982 361734
rect 20426 327818 20662 328054
rect 20746 327818 20982 328054
rect 20426 327498 20662 327734
rect 20746 327498 20982 327734
rect 20426 293818 20662 294054
rect 20746 293818 20982 294054
rect 20426 293498 20662 293734
rect 20746 293498 20982 293734
rect 20426 259818 20662 260054
rect 20746 259818 20982 260054
rect 20426 259498 20662 259734
rect 20746 259498 20982 259734
rect 20426 225818 20662 226054
rect 20746 225818 20982 226054
rect 20426 225498 20662 225734
rect 20746 225498 20982 225734
rect 20426 191818 20662 192054
rect 20746 191818 20982 192054
rect 20426 191498 20662 191734
rect 20746 191498 20982 191734
rect 20426 157818 20662 158054
rect 20746 157818 20982 158054
rect 20426 157498 20662 157734
rect 20746 157498 20982 157734
rect 20426 123818 20662 124054
rect 20746 123818 20982 124054
rect 20426 123498 20662 123734
rect 20746 123498 20982 123734
rect 20426 89818 20662 90054
rect 20746 89818 20982 90054
rect 20426 89498 20662 89734
rect 20746 89498 20982 89734
rect 20426 55818 20662 56054
rect 20746 55818 20982 56054
rect 20426 55498 20662 55734
rect 20746 55498 20982 55734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 671538 24382 671774
rect 24466 671538 24702 671774
rect 24146 671218 24382 671454
rect 24466 671218 24702 671454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 603538 24382 603774
rect 24466 603538 24702 603774
rect 24146 603218 24382 603454
rect 24466 603218 24702 603454
rect 24146 569538 24382 569774
rect 24466 569538 24702 569774
rect 24146 569218 24382 569454
rect 24466 569218 24702 569454
rect 24146 535538 24382 535774
rect 24466 535538 24702 535774
rect 24146 535218 24382 535454
rect 24466 535218 24702 535454
rect 24146 501538 24382 501774
rect 24466 501538 24702 501774
rect 24146 501218 24382 501454
rect 24466 501218 24702 501454
rect 24146 467538 24382 467774
rect 24466 467538 24702 467774
rect 24146 467218 24382 467454
rect 24466 467218 24702 467454
rect 24146 433538 24382 433774
rect 24466 433538 24702 433774
rect 24146 433218 24382 433454
rect 24466 433218 24702 433454
rect 24146 399538 24382 399774
rect 24466 399538 24702 399774
rect 24146 399218 24382 399454
rect 24466 399218 24702 399454
rect 24146 365538 24382 365774
rect 24466 365538 24702 365774
rect 24146 365218 24382 365454
rect 24466 365218 24702 365454
rect 24146 331538 24382 331774
rect 24466 331538 24702 331774
rect 24146 331218 24382 331454
rect 24466 331218 24702 331454
rect 24146 297538 24382 297774
rect 24466 297538 24702 297774
rect 24146 297218 24382 297454
rect 24466 297218 24702 297454
rect 24146 263538 24382 263774
rect 24466 263538 24702 263774
rect 24146 263218 24382 263454
rect 24466 263218 24702 263454
rect 24146 229538 24382 229774
rect 24466 229538 24702 229774
rect 24146 229218 24382 229454
rect 24466 229218 24702 229454
rect 24146 195538 24382 195774
rect 24466 195538 24702 195774
rect 24146 195218 24382 195454
rect 24466 195218 24702 195454
rect 24146 161538 24382 161774
rect 24466 161538 24702 161774
rect 24146 161218 24382 161454
rect 24466 161218 24702 161454
rect 24146 127538 24382 127774
rect 24466 127538 24702 127774
rect 24146 127218 24382 127454
rect 24466 127218 24702 127454
rect 24146 93538 24382 93774
rect 24466 93538 24702 93774
rect 24146 93218 24382 93454
rect 24466 93218 24702 93454
rect 24146 59538 24382 59774
rect 24466 59538 24702 59774
rect 24146 59218 24382 59454
rect 24466 59218 24702 59454
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 675258 28102 675494
rect 28186 675258 28422 675494
rect 27866 674938 28102 675174
rect 28186 674938 28422 675174
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 607258 28102 607494
rect 28186 607258 28422 607494
rect 27866 606938 28102 607174
rect 28186 606938 28422 607174
rect 27866 573258 28102 573494
rect 28186 573258 28422 573494
rect 27866 572938 28102 573174
rect 28186 572938 28422 573174
rect 27866 539258 28102 539494
rect 28186 539258 28422 539494
rect 27866 538938 28102 539174
rect 28186 538938 28422 539174
rect 27866 505258 28102 505494
rect 28186 505258 28422 505494
rect 27866 504938 28102 505174
rect 28186 504938 28422 505174
rect 27866 471258 28102 471494
rect 28186 471258 28422 471494
rect 27866 470938 28102 471174
rect 28186 470938 28422 471174
rect 27866 437258 28102 437494
rect 28186 437258 28422 437494
rect 27866 436938 28102 437174
rect 28186 436938 28422 437174
rect 27866 403258 28102 403494
rect 28186 403258 28422 403494
rect 27866 402938 28102 403174
rect 28186 402938 28422 403174
rect 27866 369258 28102 369494
rect 28186 369258 28422 369494
rect 27866 368938 28102 369174
rect 28186 368938 28422 369174
rect 27866 335258 28102 335494
rect 28186 335258 28422 335494
rect 27866 334938 28102 335174
rect 28186 334938 28422 335174
rect 27866 301258 28102 301494
rect 28186 301258 28422 301494
rect 27866 300938 28102 301174
rect 28186 300938 28422 301174
rect 27866 267258 28102 267494
rect 28186 267258 28422 267494
rect 27866 266938 28102 267174
rect 28186 266938 28422 267174
rect 27866 233258 28102 233494
rect 28186 233258 28422 233494
rect 27866 232938 28102 233174
rect 28186 232938 28422 233174
rect 27866 199258 28102 199494
rect 28186 199258 28422 199494
rect 27866 198938 28102 199174
rect 28186 198938 28422 199174
rect 27866 165258 28102 165494
rect 28186 165258 28422 165494
rect 27866 164938 28102 165174
rect 28186 164938 28422 165174
rect 27866 131258 28102 131494
rect 28186 131258 28422 131494
rect 27866 130938 28102 131174
rect 28186 130938 28422 131174
rect 27866 97258 28102 97494
rect 28186 97258 28422 97494
rect 27866 96938 28102 97174
rect 28186 96938 28422 97174
rect 27866 63258 28102 63494
rect 28186 63258 28422 63494
rect 27866 62938 28102 63174
rect 28186 62938 28422 63174
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 35826 704602 36062 704838
rect 36146 704602 36382 704838
rect 35826 704282 36062 704518
rect 36146 704282 36382 704518
rect 35826 683218 36062 683454
rect 36146 683218 36382 683454
rect 35826 682898 36062 683134
rect 36146 682898 36382 683134
rect 35826 649218 36062 649454
rect 36146 649218 36382 649454
rect 35826 648898 36062 649134
rect 36146 648898 36382 649134
rect 35826 615218 36062 615454
rect 36146 615218 36382 615454
rect 35826 614898 36062 615134
rect 36146 614898 36382 615134
rect 35826 581218 36062 581454
rect 36146 581218 36382 581454
rect 35826 580898 36062 581134
rect 36146 580898 36382 581134
rect 35826 547218 36062 547454
rect 36146 547218 36382 547454
rect 35826 546898 36062 547134
rect 36146 546898 36382 547134
rect 35826 513218 36062 513454
rect 36146 513218 36382 513454
rect 35826 512898 36062 513134
rect 36146 512898 36382 513134
rect 35826 479218 36062 479454
rect 36146 479218 36382 479454
rect 35826 478898 36062 479134
rect 36146 478898 36382 479134
rect 35826 445218 36062 445454
rect 36146 445218 36382 445454
rect 35826 444898 36062 445134
rect 36146 444898 36382 445134
rect 35826 411218 36062 411454
rect 36146 411218 36382 411454
rect 35826 410898 36062 411134
rect 36146 410898 36382 411134
rect 35826 377218 36062 377454
rect 36146 377218 36382 377454
rect 35826 376898 36062 377134
rect 36146 376898 36382 377134
rect 35826 343218 36062 343454
rect 36146 343218 36382 343454
rect 35826 342898 36062 343134
rect 36146 342898 36382 343134
rect 35826 309218 36062 309454
rect 36146 309218 36382 309454
rect 35826 308898 36062 309134
rect 36146 308898 36382 309134
rect 35826 275218 36062 275454
rect 36146 275218 36382 275454
rect 35826 274898 36062 275134
rect 36146 274898 36382 275134
rect 35826 241218 36062 241454
rect 36146 241218 36382 241454
rect 35826 240898 36062 241134
rect 36146 240898 36382 241134
rect 35826 207218 36062 207454
rect 36146 207218 36382 207454
rect 35826 206898 36062 207134
rect 36146 206898 36382 207134
rect 35826 173218 36062 173454
rect 36146 173218 36382 173454
rect 35826 172898 36062 173134
rect 36146 172898 36382 173134
rect 35826 139218 36062 139454
rect 36146 139218 36382 139454
rect 35826 138898 36062 139134
rect 36146 138898 36382 139134
rect 35826 105218 36062 105454
rect 36146 105218 36382 105454
rect 35826 104898 36062 105134
rect 36146 104898 36382 105134
rect 35826 71218 36062 71454
rect 36146 71218 36382 71454
rect 35826 70898 36062 71134
rect 36146 70898 36382 71134
rect 35826 37218 36062 37454
rect 36146 37218 36382 37454
rect 35826 36898 36062 37134
rect 36146 36898 36382 37134
rect 35826 3218 36062 3454
rect 36146 3218 36382 3454
rect 35826 2898 36062 3134
rect 36146 2898 36382 3134
rect 35826 -582 36062 -346
rect 36146 -582 36382 -346
rect 35826 -902 36062 -666
rect 36146 -902 36382 -666
rect 39546 705562 39782 705798
rect 39866 705562 40102 705798
rect 39546 705242 39782 705478
rect 39866 705242 40102 705478
rect 39546 686938 39782 687174
rect 39866 686938 40102 687174
rect 39546 686618 39782 686854
rect 39866 686618 40102 686854
rect 39546 652938 39782 653174
rect 39866 652938 40102 653174
rect 39546 652618 39782 652854
rect 39866 652618 40102 652854
rect 39546 618938 39782 619174
rect 39866 618938 40102 619174
rect 39546 618618 39782 618854
rect 39866 618618 40102 618854
rect 39546 584938 39782 585174
rect 39866 584938 40102 585174
rect 39546 584618 39782 584854
rect 39866 584618 40102 584854
rect 39546 550938 39782 551174
rect 39866 550938 40102 551174
rect 39546 550618 39782 550854
rect 39866 550618 40102 550854
rect 39546 516938 39782 517174
rect 39866 516938 40102 517174
rect 39546 516618 39782 516854
rect 39866 516618 40102 516854
rect 39546 482938 39782 483174
rect 39866 482938 40102 483174
rect 39546 482618 39782 482854
rect 39866 482618 40102 482854
rect 39546 448938 39782 449174
rect 39866 448938 40102 449174
rect 39546 448618 39782 448854
rect 39866 448618 40102 448854
rect 39546 414938 39782 415174
rect 39866 414938 40102 415174
rect 39546 414618 39782 414854
rect 39866 414618 40102 414854
rect 39546 380938 39782 381174
rect 39866 380938 40102 381174
rect 39546 380618 39782 380854
rect 39866 380618 40102 380854
rect 39546 346938 39782 347174
rect 39866 346938 40102 347174
rect 39546 346618 39782 346854
rect 39866 346618 40102 346854
rect 39546 312938 39782 313174
rect 39866 312938 40102 313174
rect 39546 312618 39782 312854
rect 39866 312618 40102 312854
rect 39546 278938 39782 279174
rect 39866 278938 40102 279174
rect 39546 278618 39782 278854
rect 39866 278618 40102 278854
rect 39546 244938 39782 245174
rect 39866 244938 40102 245174
rect 39546 244618 39782 244854
rect 39866 244618 40102 244854
rect 39546 210938 39782 211174
rect 39866 210938 40102 211174
rect 39546 210618 39782 210854
rect 39866 210618 40102 210854
rect 39546 176938 39782 177174
rect 39866 176938 40102 177174
rect 39546 176618 39782 176854
rect 39866 176618 40102 176854
rect 39546 142938 39782 143174
rect 39866 142938 40102 143174
rect 39546 142618 39782 142854
rect 39866 142618 40102 142854
rect 39546 108938 39782 109174
rect 39866 108938 40102 109174
rect 39546 108618 39782 108854
rect 39866 108618 40102 108854
rect 39546 74938 39782 75174
rect 39866 74938 40102 75174
rect 39546 74618 39782 74854
rect 39866 74618 40102 74854
rect 39546 40938 39782 41174
rect 39866 40938 40102 41174
rect 39546 40618 39782 40854
rect 39866 40618 40102 40854
rect 39546 6938 39782 7174
rect 39866 6938 40102 7174
rect 39546 6618 39782 6854
rect 39866 6618 40102 6854
rect 39546 -1542 39782 -1306
rect 39866 -1542 40102 -1306
rect 39546 -1862 39782 -1626
rect 39866 -1862 40102 -1626
rect 43266 706522 43502 706758
rect 43586 706522 43822 706758
rect 43266 706202 43502 706438
rect 43586 706202 43822 706438
rect 43266 690658 43502 690894
rect 43586 690658 43822 690894
rect 43266 690338 43502 690574
rect 43586 690338 43822 690574
rect 43266 656658 43502 656894
rect 43586 656658 43822 656894
rect 43266 656338 43502 656574
rect 43586 656338 43822 656574
rect 43266 622658 43502 622894
rect 43586 622658 43822 622894
rect 43266 622338 43502 622574
rect 43586 622338 43822 622574
rect 43266 588658 43502 588894
rect 43586 588658 43822 588894
rect 43266 588338 43502 588574
rect 43586 588338 43822 588574
rect 43266 554658 43502 554894
rect 43586 554658 43822 554894
rect 43266 554338 43502 554574
rect 43586 554338 43822 554574
rect 43266 520658 43502 520894
rect 43586 520658 43822 520894
rect 43266 520338 43502 520574
rect 43586 520338 43822 520574
rect 43266 486658 43502 486894
rect 43586 486658 43822 486894
rect 43266 486338 43502 486574
rect 43586 486338 43822 486574
rect 43266 452658 43502 452894
rect 43586 452658 43822 452894
rect 43266 452338 43502 452574
rect 43586 452338 43822 452574
rect 43266 418658 43502 418894
rect 43586 418658 43822 418894
rect 43266 418338 43502 418574
rect 43586 418338 43822 418574
rect 43266 384658 43502 384894
rect 43586 384658 43822 384894
rect 43266 384338 43502 384574
rect 43586 384338 43822 384574
rect 43266 350658 43502 350894
rect 43586 350658 43822 350894
rect 43266 350338 43502 350574
rect 43586 350338 43822 350574
rect 43266 316658 43502 316894
rect 43586 316658 43822 316894
rect 43266 316338 43502 316574
rect 43586 316338 43822 316574
rect 43266 282658 43502 282894
rect 43586 282658 43822 282894
rect 43266 282338 43502 282574
rect 43586 282338 43822 282574
rect 43266 248658 43502 248894
rect 43586 248658 43822 248894
rect 43266 248338 43502 248574
rect 43586 248338 43822 248574
rect 46986 707482 47222 707718
rect 47306 707482 47542 707718
rect 46986 707162 47222 707398
rect 47306 707162 47542 707398
rect 46986 694378 47222 694614
rect 47306 694378 47542 694614
rect 46986 694058 47222 694294
rect 47306 694058 47542 694294
rect 46986 660378 47222 660614
rect 47306 660378 47542 660614
rect 46986 660058 47222 660294
rect 47306 660058 47542 660294
rect 46986 626378 47222 626614
rect 47306 626378 47542 626614
rect 46986 626058 47222 626294
rect 47306 626058 47542 626294
rect 46986 592378 47222 592614
rect 47306 592378 47542 592614
rect 46986 592058 47222 592294
rect 47306 592058 47542 592294
rect 46986 558378 47222 558614
rect 47306 558378 47542 558614
rect 46986 558058 47222 558294
rect 47306 558058 47542 558294
rect 46986 524378 47222 524614
rect 47306 524378 47542 524614
rect 46986 524058 47222 524294
rect 47306 524058 47542 524294
rect 46986 490378 47222 490614
rect 47306 490378 47542 490614
rect 46986 490058 47222 490294
rect 47306 490058 47542 490294
rect 46986 456378 47222 456614
rect 47306 456378 47542 456614
rect 46986 456058 47222 456294
rect 47306 456058 47542 456294
rect 46986 422378 47222 422614
rect 47306 422378 47542 422614
rect 46986 422058 47222 422294
rect 47306 422058 47542 422294
rect 46986 388378 47222 388614
rect 47306 388378 47542 388614
rect 46986 388058 47222 388294
rect 47306 388058 47542 388294
rect 46986 354378 47222 354614
rect 47306 354378 47542 354614
rect 46986 354058 47222 354294
rect 47306 354058 47542 354294
rect 46986 320378 47222 320614
rect 47306 320378 47542 320614
rect 46986 320058 47222 320294
rect 47306 320058 47542 320294
rect 46986 286378 47222 286614
rect 47306 286378 47542 286614
rect 46986 286058 47222 286294
rect 47306 286058 47542 286294
rect 46986 252378 47222 252614
rect 47306 252378 47542 252614
rect 46986 252058 47222 252294
rect 47306 252058 47542 252294
rect 50706 708442 50942 708678
rect 51026 708442 51262 708678
rect 50706 708122 50942 708358
rect 51026 708122 51262 708358
rect 50706 698098 50942 698334
rect 51026 698098 51262 698334
rect 50706 697778 50942 698014
rect 51026 697778 51262 698014
rect 50706 664098 50942 664334
rect 51026 664098 51262 664334
rect 50706 663778 50942 664014
rect 51026 663778 51262 664014
rect 50706 630098 50942 630334
rect 51026 630098 51262 630334
rect 50706 629778 50942 630014
rect 51026 629778 51262 630014
rect 50706 596098 50942 596334
rect 51026 596098 51262 596334
rect 50706 595778 50942 596014
rect 51026 595778 51262 596014
rect 50706 562098 50942 562334
rect 51026 562098 51262 562334
rect 50706 561778 50942 562014
rect 51026 561778 51262 562014
rect 50706 528098 50942 528334
rect 51026 528098 51262 528334
rect 50706 527778 50942 528014
rect 51026 527778 51262 528014
rect 50706 494098 50942 494334
rect 51026 494098 51262 494334
rect 50706 493778 50942 494014
rect 51026 493778 51262 494014
rect 50706 460098 50942 460334
rect 51026 460098 51262 460334
rect 50706 459778 50942 460014
rect 51026 459778 51262 460014
rect 50706 426098 50942 426334
rect 51026 426098 51262 426334
rect 50706 425778 50942 426014
rect 51026 425778 51262 426014
rect 50706 392098 50942 392334
rect 51026 392098 51262 392334
rect 50706 391778 50942 392014
rect 51026 391778 51262 392014
rect 50706 358098 50942 358334
rect 51026 358098 51262 358334
rect 50706 357778 50942 358014
rect 51026 357778 51262 358014
rect 50706 324098 50942 324334
rect 51026 324098 51262 324334
rect 50706 323778 50942 324014
rect 51026 323778 51262 324014
rect 50706 290098 50942 290334
rect 51026 290098 51262 290334
rect 50706 289778 50942 290014
rect 51026 289778 51262 290014
rect 50706 256098 50942 256334
rect 51026 256098 51262 256334
rect 50706 255778 50942 256014
rect 51026 255778 51262 256014
rect 54426 709402 54662 709638
rect 54746 709402 54982 709638
rect 54426 709082 54662 709318
rect 54746 709082 54982 709318
rect 54426 667818 54662 668054
rect 54746 667818 54982 668054
rect 54426 667498 54662 667734
rect 54746 667498 54982 667734
rect 54426 633818 54662 634054
rect 54746 633818 54982 634054
rect 54426 633498 54662 633734
rect 54746 633498 54982 633734
rect 54426 599818 54662 600054
rect 54746 599818 54982 600054
rect 54426 599498 54662 599734
rect 54746 599498 54982 599734
rect 54426 565818 54662 566054
rect 54746 565818 54982 566054
rect 54426 565498 54662 565734
rect 54746 565498 54982 565734
rect 54426 531818 54662 532054
rect 54746 531818 54982 532054
rect 54426 531498 54662 531734
rect 54746 531498 54982 531734
rect 54426 497818 54662 498054
rect 54746 497818 54982 498054
rect 54426 497498 54662 497734
rect 54746 497498 54982 497734
rect 54426 463818 54662 464054
rect 54746 463818 54982 464054
rect 54426 463498 54662 463734
rect 54746 463498 54982 463734
rect 54426 429818 54662 430054
rect 54746 429818 54982 430054
rect 54426 429498 54662 429734
rect 54746 429498 54982 429734
rect 54426 395818 54662 396054
rect 54746 395818 54982 396054
rect 54426 395498 54662 395734
rect 54746 395498 54982 395734
rect 54426 361818 54662 362054
rect 54746 361818 54982 362054
rect 54426 361498 54662 361734
rect 54746 361498 54982 361734
rect 54426 327818 54662 328054
rect 54746 327818 54982 328054
rect 54426 327498 54662 327734
rect 54746 327498 54982 327734
rect 54426 293818 54662 294054
rect 54746 293818 54982 294054
rect 54426 293498 54662 293734
rect 54746 293498 54982 293734
rect 54426 259818 54662 260054
rect 54746 259818 54982 260054
rect 54426 259498 54662 259734
rect 54746 259498 54982 259734
rect 54426 225705 54662 225941
rect 54746 225705 54982 225941
rect 58146 710362 58382 710598
rect 58466 710362 58702 710598
rect 58146 710042 58382 710278
rect 58466 710042 58702 710278
rect 58146 671538 58382 671774
rect 58466 671538 58702 671774
rect 58146 671218 58382 671454
rect 58466 671218 58702 671454
rect 58146 637538 58382 637774
rect 58466 637538 58702 637774
rect 58146 637218 58382 637454
rect 58466 637218 58702 637454
rect 58146 603538 58382 603774
rect 58466 603538 58702 603774
rect 58146 603218 58382 603454
rect 58466 603218 58702 603454
rect 58146 569538 58382 569774
rect 58466 569538 58702 569774
rect 58146 569218 58382 569454
rect 58466 569218 58702 569454
rect 58146 535538 58382 535774
rect 58466 535538 58702 535774
rect 58146 535218 58382 535454
rect 58466 535218 58702 535454
rect 58146 501538 58382 501774
rect 58466 501538 58702 501774
rect 58146 501218 58382 501454
rect 58466 501218 58702 501454
rect 58146 467538 58382 467774
rect 58466 467538 58702 467774
rect 58146 467218 58382 467454
rect 58466 467218 58702 467454
rect 58146 433538 58382 433774
rect 58466 433538 58702 433774
rect 58146 433218 58382 433454
rect 58466 433218 58702 433454
rect 58146 399538 58382 399774
rect 58466 399538 58702 399774
rect 58146 399218 58382 399454
rect 58466 399218 58702 399454
rect 58146 365538 58382 365774
rect 58466 365538 58702 365774
rect 58146 365218 58382 365454
rect 58466 365218 58702 365454
rect 58146 331538 58382 331774
rect 58466 331538 58702 331774
rect 58146 331218 58382 331454
rect 58466 331218 58702 331454
rect 58146 297538 58382 297774
rect 58466 297538 58702 297774
rect 58146 297218 58382 297454
rect 58466 297218 58702 297454
rect 58146 263538 58382 263774
rect 58466 263538 58702 263774
rect 58146 263218 58382 263454
rect 58466 263218 58702 263454
rect 58146 229538 58382 229774
rect 58466 229538 58702 229774
rect 58146 229218 58382 229454
rect 58466 229218 58702 229454
rect 61866 711322 62102 711558
rect 62186 711322 62422 711558
rect 61866 711002 62102 711238
rect 62186 711002 62422 711238
rect 61866 675258 62102 675494
rect 62186 675258 62422 675494
rect 61866 674938 62102 675174
rect 62186 674938 62422 675174
rect 61866 641258 62102 641494
rect 62186 641258 62422 641494
rect 61866 640938 62102 641174
rect 62186 640938 62422 641174
rect 61866 607258 62102 607494
rect 62186 607258 62422 607494
rect 61866 606938 62102 607174
rect 62186 606938 62422 607174
rect 61866 573258 62102 573494
rect 62186 573258 62422 573494
rect 61866 572938 62102 573174
rect 62186 572938 62422 573174
rect 61866 539258 62102 539494
rect 62186 539258 62422 539494
rect 61866 538938 62102 539174
rect 62186 538938 62422 539174
rect 61866 505258 62102 505494
rect 62186 505258 62422 505494
rect 61866 504938 62102 505174
rect 62186 504938 62422 505174
rect 61866 471258 62102 471494
rect 62186 471258 62422 471494
rect 61866 470938 62102 471174
rect 62186 470938 62422 471174
rect 61866 437258 62102 437494
rect 62186 437258 62422 437494
rect 61866 436938 62102 437174
rect 62186 436938 62422 437174
rect 61866 403258 62102 403494
rect 62186 403258 62422 403494
rect 61866 402938 62102 403174
rect 62186 402938 62422 403174
rect 61866 369258 62102 369494
rect 62186 369258 62422 369494
rect 61866 368938 62102 369174
rect 62186 368938 62422 369174
rect 61866 335258 62102 335494
rect 62186 335258 62422 335494
rect 61866 334938 62102 335174
rect 62186 334938 62422 335174
rect 61866 301258 62102 301494
rect 62186 301258 62422 301494
rect 61866 300938 62102 301174
rect 62186 300938 62422 301174
rect 61866 267258 62102 267494
rect 62186 267258 62422 267494
rect 61866 266938 62102 267174
rect 62186 266938 62422 267174
rect 61866 233258 62102 233494
rect 62186 233258 62422 233494
rect 61866 232938 62102 233174
rect 62186 232938 62422 233174
rect 69826 704602 70062 704838
rect 70146 704602 70382 704838
rect 69826 704282 70062 704518
rect 70146 704282 70382 704518
rect 69826 683218 70062 683454
rect 70146 683218 70382 683454
rect 69826 682898 70062 683134
rect 70146 682898 70382 683134
rect 69826 649218 70062 649454
rect 70146 649218 70382 649454
rect 69826 648898 70062 649134
rect 70146 648898 70382 649134
rect 69826 615218 70062 615454
rect 70146 615218 70382 615454
rect 69826 614898 70062 615134
rect 70146 614898 70382 615134
rect 69826 581218 70062 581454
rect 70146 581218 70382 581454
rect 69826 580898 70062 581134
rect 70146 580898 70382 581134
rect 69826 547218 70062 547454
rect 70146 547218 70382 547454
rect 69826 546898 70062 547134
rect 70146 546898 70382 547134
rect 69826 513218 70062 513454
rect 70146 513218 70382 513454
rect 69826 512898 70062 513134
rect 70146 512898 70382 513134
rect 69826 479218 70062 479454
rect 70146 479218 70382 479454
rect 69826 478898 70062 479134
rect 70146 478898 70382 479134
rect 69826 445218 70062 445454
rect 70146 445218 70382 445454
rect 69826 444898 70062 445134
rect 70146 444898 70382 445134
rect 69826 411218 70062 411454
rect 70146 411218 70382 411454
rect 69826 410898 70062 411134
rect 70146 410898 70382 411134
rect 69826 377218 70062 377454
rect 70146 377218 70382 377454
rect 69826 376898 70062 377134
rect 70146 376898 70382 377134
rect 69826 343218 70062 343454
rect 70146 343218 70382 343454
rect 69826 342898 70062 343134
rect 70146 342898 70382 343134
rect 69826 309218 70062 309454
rect 70146 309218 70382 309454
rect 69826 308898 70062 309134
rect 70146 308898 70382 309134
rect 69826 275218 70062 275454
rect 70146 275218 70382 275454
rect 69826 274898 70062 275134
rect 70146 274898 70382 275134
rect 69826 241218 70062 241454
rect 70146 241218 70382 241454
rect 69826 240898 70062 241134
rect 70146 240898 70382 241134
rect 73546 705562 73782 705798
rect 73866 705562 74102 705798
rect 73546 705242 73782 705478
rect 73866 705242 74102 705478
rect 73546 686938 73782 687174
rect 73866 686938 74102 687174
rect 73546 686618 73782 686854
rect 73866 686618 74102 686854
rect 73546 652938 73782 653174
rect 73866 652938 74102 653174
rect 73546 652618 73782 652854
rect 73866 652618 74102 652854
rect 73546 618938 73782 619174
rect 73866 618938 74102 619174
rect 73546 618618 73782 618854
rect 73866 618618 74102 618854
rect 73546 584938 73782 585174
rect 73866 584938 74102 585174
rect 73546 584618 73782 584854
rect 73866 584618 74102 584854
rect 73546 550938 73782 551174
rect 73866 550938 74102 551174
rect 73546 550618 73782 550854
rect 73866 550618 74102 550854
rect 73546 516938 73782 517174
rect 73866 516938 74102 517174
rect 73546 516618 73782 516854
rect 73866 516618 74102 516854
rect 73546 482938 73782 483174
rect 73866 482938 74102 483174
rect 73546 482618 73782 482854
rect 73866 482618 74102 482854
rect 73546 448938 73782 449174
rect 73866 448938 74102 449174
rect 73546 448618 73782 448854
rect 73866 448618 74102 448854
rect 73546 414938 73782 415174
rect 73866 414938 74102 415174
rect 73546 414618 73782 414854
rect 73866 414618 74102 414854
rect 73546 380938 73782 381174
rect 73866 380938 74102 381174
rect 73546 380618 73782 380854
rect 73866 380618 74102 380854
rect 73546 346938 73782 347174
rect 73866 346938 74102 347174
rect 73546 346618 73782 346854
rect 73866 346618 74102 346854
rect 73546 312938 73782 313174
rect 73866 312938 74102 313174
rect 73546 312618 73782 312854
rect 73866 312618 74102 312854
rect 73546 278938 73782 279174
rect 73866 278938 74102 279174
rect 73546 278618 73782 278854
rect 73866 278618 74102 278854
rect 73546 244938 73782 245174
rect 73866 244938 74102 245174
rect 73546 244618 73782 244854
rect 73866 244618 74102 244854
rect 65339 229535 65575 229771
rect 65659 229535 65895 229771
rect 65979 229535 66215 229771
rect 66299 229535 66535 229771
rect 66619 229535 66855 229771
rect 66939 229535 67175 229771
rect 67259 229535 67495 229771
rect 67579 229535 67815 229771
rect 67899 229535 68135 229771
rect 68219 229535 68455 229771
rect 68539 229535 68775 229771
rect 68859 229535 69095 229771
rect 69179 229535 69415 229771
rect 69499 229535 69735 229771
rect 69819 229535 70055 229771
rect 65339 229215 65575 229451
rect 65659 229215 65895 229451
rect 65979 229215 66215 229451
rect 66299 229215 66535 229451
rect 66619 229215 66855 229451
rect 66939 229215 67175 229451
rect 67259 229215 67495 229451
rect 67579 229215 67815 229451
rect 67899 229215 68135 229451
rect 68219 229215 68455 229451
rect 68539 229215 68775 229451
rect 68859 229215 69095 229451
rect 69179 229215 69415 229451
rect 69499 229215 69735 229451
rect 69819 229215 70055 229451
rect 65462 225565 65698 225801
rect 65782 225565 66018 225801
rect 66102 225565 66338 225801
rect 66422 225565 66658 225801
rect 66742 225565 66978 225801
rect 67062 225565 67298 225801
rect 67382 225565 67618 225801
rect 67702 225565 67938 225801
rect 68022 225565 68258 225801
rect 68342 225565 68578 225801
rect 68662 225565 68898 225801
rect 68982 225565 69218 225801
rect 69302 225565 69538 225801
rect 69622 225565 69858 225801
rect 69942 225565 70178 225801
rect 70262 225565 70498 225801
rect 70582 225565 70818 225801
rect 70902 225565 71138 225801
rect 77266 706522 77502 706758
rect 77586 706522 77822 706758
rect 77266 706202 77502 706438
rect 77586 706202 77822 706438
rect 77266 690658 77502 690894
rect 77586 690658 77822 690894
rect 77266 690338 77502 690574
rect 77586 690338 77822 690574
rect 77266 656658 77502 656894
rect 77586 656658 77822 656894
rect 77266 656338 77502 656574
rect 77586 656338 77822 656574
rect 77266 622658 77502 622894
rect 77586 622658 77822 622894
rect 77266 622338 77502 622574
rect 77586 622338 77822 622574
rect 77266 588658 77502 588894
rect 77586 588658 77822 588894
rect 77266 588338 77502 588574
rect 77586 588338 77822 588574
rect 77266 554658 77502 554894
rect 77586 554658 77822 554894
rect 77266 554338 77502 554574
rect 77586 554338 77822 554574
rect 77266 520658 77502 520894
rect 77586 520658 77822 520894
rect 77266 520338 77502 520574
rect 77586 520338 77822 520574
rect 77266 486658 77502 486894
rect 77586 486658 77822 486894
rect 77266 486338 77502 486574
rect 77586 486338 77822 486574
rect 77266 452658 77502 452894
rect 77586 452658 77822 452894
rect 77266 452338 77502 452574
rect 77586 452338 77822 452574
rect 77266 418658 77502 418894
rect 77586 418658 77822 418894
rect 77266 418338 77502 418574
rect 77586 418338 77822 418574
rect 77266 384658 77502 384894
rect 77586 384658 77822 384894
rect 77266 384338 77502 384574
rect 77586 384338 77822 384574
rect 77266 350658 77502 350894
rect 77586 350658 77822 350894
rect 77266 350338 77502 350574
rect 77586 350338 77822 350574
rect 77266 316658 77502 316894
rect 77586 316658 77822 316894
rect 77266 316338 77502 316574
rect 77586 316338 77822 316574
rect 77266 282658 77502 282894
rect 77586 282658 77822 282894
rect 77266 282338 77502 282574
rect 77586 282338 77822 282574
rect 77266 248658 77502 248894
rect 77586 248658 77822 248894
rect 77266 248338 77502 248574
rect 77586 248338 77822 248574
rect 80986 707482 81222 707718
rect 81306 707482 81542 707718
rect 80986 707162 81222 707398
rect 81306 707162 81542 707398
rect 80986 694378 81222 694614
rect 81306 694378 81542 694614
rect 80986 694058 81222 694294
rect 81306 694058 81542 694294
rect 80986 660378 81222 660614
rect 81306 660378 81542 660614
rect 80986 660058 81222 660294
rect 81306 660058 81542 660294
rect 80986 626378 81222 626614
rect 81306 626378 81542 626614
rect 80986 626058 81222 626294
rect 81306 626058 81542 626294
rect 80986 592378 81222 592614
rect 81306 592378 81542 592614
rect 80986 592058 81222 592294
rect 81306 592058 81542 592294
rect 80986 558378 81222 558614
rect 81306 558378 81542 558614
rect 80986 558058 81222 558294
rect 81306 558058 81542 558294
rect 80986 524378 81222 524614
rect 81306 524378 81542 524614
rect 80986 524058 81222 524294
rect 81306 524058 81542 524294
rect 80986 490378 81222 490614
rect 81306 490378 81542 490614
rect 80986 490058 81222 490294
rect 81306 490058 81542 490294
rect 80986 456378 81222 456614
rect 81306 456378 81542 456614
rect 80986 456058 81222 456294
rect 81306 456058 81542 456294
rect 80986 422378 81222 422614
rect 81306 422378 81542 422614
rect 80986 422058 81222 422294
rect 81306 422058 81542 422294
rect 80986 388378 81222 388614
rect 81306 388378 81542 388614
rect 80986 388058 81222 388294
rect 81306 388058 81542 388294
rect 80986 354378 81222 354614
rect 81306 354378 81542 354614
rect 80986 354058 81222 354294
rect 81306 354058 81542 354294
rect 80986 320378 81222 320614
rect 81306 320378 81542 320614
rect 80986 320058 81222 320294
rect 81306 320058 81542 320294
rect 80986 286378 81222 286614
rect 81306 286378 81542 286614
rect 80986 286058 81222 286294
rect 81306 286058 81542 286294
rect 80986 252378 81222 252614
rect 81306 252378 81542 252614
rect 80986 252058 81222 252294
rect 81306 252058 81542 252294
rect 84706 708442 84942 708678
rect 85026 708442 85262 708678
rect 84706 708122 84942 708358
rect 85026 708122 85262 708358
rect 84706 698098 84942 698334
rect 85026 698098 85262 698334
rect 84706 697778 84942 698014
rect 85026 697778 85262 698014
rect 84706 664098 84942 664334
rect 85026 664098 85262 664334
rect 84706 663778 84942 664014
rect 85026 663778 85262 664014
rect 84706 630098 84942 630334
rect 85026 630098 85262 630334
rect 84706 629778 84942 630014
rect 85026 629778 85262 630014
rect 84706 596098 84942 596334
rect 85026 596098 85262 596334
rect 84706 595778 84942 596014
rect 85026 595778 85262 596014
rect 84706 562098 84942 562334
rect 85026 562098 85262 562334
rect 84706 561778 84942 562014
rect 85026 561778 85262 562014
rect 84706 528098 84942 528334
rect 85026 528098 85262 528334
rect 84706 527778 84942 528014
rect 85026 527778 85262 528014
rect 84706 494098 84942 494334
rect 85026 494098 85262 494334
rect 84706 493778 84942 494014
rect 85026 493778 85262 494014
rect 84706 460098 84942 460334
rect 85026 460098 85262 460334
rect 84706 459778 84942 460014
rect 85026 459778 85262 460014
rect 84706 426098 84942 426334
rect 85026 426098 85262 426334
rect 84706 425778 84942 426014
rect 85026 425778 85262 426014
rect 84706 392098 84942 392334
rect 85026 392098 85262 392334
rect 84706 391778 84942 392014
rect 85026 391778 85262 392014
rect 84706 358098 84942 358334
rect 85026 358098 85262 358334
rect 84706 357778 84942 358014
rect 85026 357778 85262 358014
rect 84706 324098 84942 324334
rect 85026 324098 85262 324334
rect 84706 323778 84942 324014
rect 85026 323778 85262 324014
rect 84706 290098 84942 290334
rect 85026 290098 85262 290334
rect 84706 289778 84942 290014
rect 85026 289778 85262 290014
rect 84706 256098 84942 256334
rect 85026 256098 85262 256334
rect 84706 255778 84942 256014
rect 85026 255778 85262 256014
rect 88426 709402 88662 709638
rect 88746 709402 88982 709638
rect 88426 709082 88662 709318
rect 88746 709082 88982 709318
rect 88426 667818 88662 668054
rect 88746 667818 88982 668054
rect 88426 667498 88662 667734
rect 88746 667498 88982 667734
rect 88426 633818 88662 634054
rect 88746 633818 88982 634054
rect 88426 633498 88662 633734
rect 88746 633498 88982 633734
rect 88426 599818 88662 600054
rect 88746 599818 88982 600054
rect 88426 599498 88662 599734
rect 88746 599498 88982 599734
rect 88426 565818 88662 566054
rect 88746 565818 88982 566054
rect 88426 565498 88662 565734
rect 88746 565498 88982 565734
rect 88426 531818 88662 532054
rect 88746 531818 88982 532054
rect 88426 531498 88662 531734
rect 88746 531498 88982 531734
rect 88426 497818 88662 498054
rect 88746 497818 88982 498054
rect 88426 497498 88662 497734
rect 88746 497498 88982 497734
rect 88426 463818 88662 464054
rect 88746 463818 88982 464054
rect 88426 463498 88662 463734
rect 88746 463498 88982 463734
rect 88426 429818 88662 430054
rect 88746 429818 88982 430054
rect 88426 429498 88662 429734
rect 88746 429498 88982 429734
rect 88426 395818 88662 396054
rect 88746 395818 88982 396054
rect 88426 395498 88662 395734
rect 88746 395498 88982 395734
rect 88426 361818 88662 362054
rect 88746 361818 88982 362054
rect 88426 361498 88662 361734
rect 88746 361498 88982 361734
rect 88426 327818 88662 328054
rect 88746 327818 88982 328054
rect 88426 327498 88662 327734
rect 88746 327498 88982 327734
rect 88426 293818 88662 294054
rect 88746 293818 88982 294054
rect 88426 293498 88662 293734
rect 88746 293498 88982 293734
rect 88426 259818 88662 260054
rect 88746 259818 88982 260054
rect 88426 259498 88662 259734
rect 88746 259498 88982 259734
rect 88426 225755 88662 225991
rect 88746 225755 88982 225991
rect 92146 710362 92382 710598
rect 92466 710362 92702 710598
rect 92146 710042 92382 710278
rect 92466 710042 92702 710278
rect 92146 671538 92382 671774
rect 92466 671538 92702 671774
rect 92146 671218 92382 671454
rect 92466 671218 92702 671454
rect 92146 637538 92382 637774
rect 92466 637538 92702 637774
rect 92146 637218 92382 637454
rect 92466 637218 92702 637454
rect 92146 603538 92382 603774
rect 92466 603538 92702 603774
rect 92146 603218 92382 603454
rect 92466 603218 92702 603454
rect 92146 569538 92382 569774
rect 92466 569538 92702 569774
rect 92146 569218 92382 569454
rect 92466 569218 92702 569454
rect 92146 535538 92382 535774
rect 92466 535538 92702 535774
rect 92146 535218 92382 535454
rect 92466 535218 92702 535454
rect 92146 501538 92382 501774
rect 92466 501538 92702 501774
rect 92146 501218 92382 501454
rect 92466 501218 92702 501454
rect 92146 467538 92382 467774
rect 92466 467538 92702 467774
rect 92146 467218 92382 467454
rect 92466 467218 92702 467454
rect 92146 433538 92382 433774
rect 92466 433538 92702 433774
rect 92146 433218 92382 433454
rect 92466 433218 92702 433454
rect 92146 399538 92382 399774
rect 92466 399538 92702 399774
rect 92146 399218 92382 399454
rect 92466 399218 92702 399454
rect 92146 365538 92382 365774
rect 92466 365538 92702 365774
rect 92146 365218 92382 365454
rect 92466 365218 92702 365454
rect 92146 331538 92382 331774
rect 92466 331538 92702 331774
rect 92146 331218 92382 331454
rect 92466 331218 92702 331454
rect 92146 297538 92382 297774
rect 92466 297538 92702 297774
rect 92146 297218 92382 297454
rect 92466 297218 92702 297454
rect 92146 263538 92382 263774
rect 92466 263538 92702 263774
rect 92146 263218 92382 263454
rect 92466 263218 92702 263454
rect 92146 229538 92382 229774
rect 92466 229538 92702 229774
rect 92146 229218 92382 229454
rect 92466 229218 92702 229454
rect 95866 711322 96102 711558
rect 96186 711322 96422 711558
rect 95866 711002 96102 711238
rect 96186 711002 96422 711238
rect 95866 675258 96102 675494
rect 96186 675258 96422 675494
rect 95866 674938 96102 675174
rect 96186 674938 96422 675174
rect 95866 641258 96102 641494
rect 96186 641258 96422 641494
rect 95866 640938 96102 641174
rect 96186 640938 96422 641174
rect 95866 607258 96102 607494
rect 96186 607258 96422 607494
rect 95866 606938 96102 607174
rect 96186 606938 96422 607174
rect 95866 573258 96102 573494
rect 96186 573258 96422 573494
rect 95866 572938 96102 573174
rect 96186 572938 96422 573174
rect 95866 539258 96102 539494
rect 96186 539258 96422 539494
rect 95866 538938 96102 539174
rect 96186 538938 96422 539174
rect 95866 505258 96102 505494
rect 96186 505258 96422 505494
rect 95866 504938 96102 505174
rect 96186 504938 96422 505174
rect 95866 471258 96102 471494
rect 96186 471258 96422 471494
rect 95866 470938 96102 471174
rect 96186 470938 96422 471174
rect 95866 437258 96102 437494
rect 96186 437258 96422 437494
rect 95866 436938 96102 437174
rect 96186 436938 96422 437174
rect 95866 403258 96102 403494
rect 96186 403258 96422 403494
rect 95866 402938 96102 403174
rect 96186 402938 96422 403174
rect 95866 369258 96102 369494
rect 96186 369258 96422 369494
rect 95866 368938 96102 369174
rect 96186 368938 96422 369174
rect 95866 335258 96102 335494
rect 96186 335258 96422 335494
rect 95866 334938 96102 335174
rect 96186 334938 96422 335174
rect 95866 301258 96102 301494
rect 96186 301258 96422 301494
rect 95866 300938 96102 301174
rect 96186 300938 96422 301174
rect 95866 267258 96102 267494
rect 96186 267258 96422 267494
rect 95866 266938 96102 267174
rect 96186 266938 96422 267174
rect 95866 233258 96102 233494
rect 96186 233258 96422 233494
rect 95866 232938 96102 233174
rect 96186 232938 96422 233174
rect 103826 704602 104062 704838
rect 104146 704602 104382 704838
rect 103826 704282 104062 704518
rect 104146 704282 104382 704518
rect 103826 683218 104062 683454
rect 104146 683218 104382 683454
rect 103826 682898 104062 683134
rect 104146 682898 104382 683134
rect 103826 649218 104062 649454
rect 104146 649218 104382 649454
rect 103826 648898 104062 649134
rect 104146 648898 104382 649134
rect 103826 615218 104062 615454
rect 104146 615218 104382 615454
rect 103826 614898 104062 615134
rect 104146 614898 104382 615134
rect 103826 581218 104062 581454
rect 104146 581218 104382 581454
rect 103826 580898 104062 581134
rect 104146 580898 104382 581134
rect 103826 547218 104062 547454
rect 104146 547218 104382 547454
rect 103826 546898 104062 547134
rect 104146 546898 104382 547134
rect 103826 513218 104062 513454
rect 104146 513218 104382 513454
rect 103826 512898 104062 513134
rect 104146 512898 104382 513134
rect 103826 479218 104062 479454
rect 104146 479218 104382 479454
rect 103826 478898 104062 479134
rect 104146 478898 104382 479134
rect 103826 445218 104062 445454
rect 104146 445218 104382 445454
rect 103826 444898 104062 445134
rect 104146 444898 104382 445134
rect 103826 411218 104062 411454
rect 104146 411218 104382 411454
rect 103826 410898 104062 411134
rect 104146 410898 104382 411134
rect 103826 377218 104062 377454
rect 104146 377218 104382 377454
rect 103826 376898 104062 377134
rect 104146 376898 104382 377134
rect 103826 343218 104062 343454
rect 104146 343218 104382 343454
rect 103826 342898 104062 343134
rect 104146 342898 104382 343134
rect 103826 309218 104062 309454
rect 104146 309218 104382 309454
rect 103826 308898 104062 309134
rect 104146 308898 104382 309134
rect 103826 275218 104062 275454
rect 104146 275218 104382 275454
rect 103826 274898 104062 275134
rect 104146 274898 104382 275134
rect 103826 241218 104062 241454
rect 104146 241218 104382 241454
rect 103826 240898 104062 241134
rect 104146 240898 104382 241134
rect 107546 705562 107782 705798
rect 107866 705562 108102 705798
rect 107546 705242 107782 705478
rect 107866 705242 108102 705478
rect 107546 686938 107782 687174
rect 107866 686938 108102 687174
rect 107546 686618 107782 686854
rect 107866 686618 108102 686854
rect 107546 652938 107782 653174
rect 107866 652938 108102 653174
rect 107546 652618 107782 652854
rect 107866 652618 108102 652854
rect 107546 618938 107782 619174
rect 107866 618938 108102 619174
rect 107546 618618 107782 618854
rect 107866 618618 108102 618854
rect 107546 584938 107782 585174
rect 107866 584938 108102 585174
rect 107546 584618 107782 584854
rect 107866 584618 108102 584854
rect 107546 550938 107782 551174
rect 107866 550938 108102 551174
rect 107546 550618 107782 550854
rect 107866 550618 108102 550854
rect 107546 516938 107782 517174
rect 107866 516938 108102 517174
rect 107546 516618 107782 516854
rect 107866 516618 108102 516854
rect 107546 482938 107782 483174
rect 107866 482938 108102 483174
rect 107546 482618 107782 482854
rect 107866 482618 108102 482854
rect 107546 448938 107782 449174
rect 107866 448938 108102 449174
rect 107546 448618 107782 448854
rect 107866 448618 108102 448854
rect 107546 414938 107782 415174
rect 107866 414938 108102 415174
rect 107546 414618 107782 414854
rect 107866 414618 108102 414854
rect 107546 380938 107782 381174
rect 107866 380938 108102 381174
rect 107546 380618 107782 380854
rect 107866 380618 108102 380854
rect 107546 346938 107782 347174
rect 107866 346938 108102 347174
rect 107546 346618 107782 346854
rect 107866 346618 108102 346854
rect 107546 312938 107782 313174
rect 107866 312938 108102 313174
rect 107546 312618 107782 312854
rect 107866 312618 108102 312854
rect 107546 278938 107782 279174
rect 107866 278938 108102 279174
rect 107546 278618 107782 278854
rect 107866 278618 108102 278854
rect 107546 244938 107782 245174
rect 107866 244938 108102 245174
rect 107546 244618 107782 244854
rect 107866 244618 108102 244854
rect 111266 706522 111502 706758
rect 111586 706522 111822 706758
rect 111266 706202 111502 706438
rect 111586 706202 111822 706438
rect 111266 690658 111502 690894
rect 111586 690658 111822 690894
rect 111266 690338 111502 690574
rect 111586 690338 111822 690574
rect 111266 656658 111502 656894
rect 111586 656658 111822 656894
rect 111266 656338 111502 656574
rect 111586 656338 111822 656574
rect 111266 622658 111502 622894
rect 111586 622658 111822 622894
rect 111266 622338 111502 622574
rect 111586 622338 111822 622574
rect 111266 588658 111502 588894
rect 111586 588658 111822 588894
rect 111266 588338 111502 588574
rect 111586 588338 111822 588574
rect 111266 554658 111502 554894
rect 111586 554658 111822 554894
rect 111266 554338 111502 554574
rect 111586 554338 111822 554574
rect 111266 520658 111502 520894
rect 111586 520658 111822 520894
rect 111266 520338 111502 520574
rect 111586 520338 111822 520574
rect 111266 486658 111502 486894
rect 111586 486658 111822 486894
rect 111266 486338 111502 486574
rect 111586 486338 111822 486574
rect 111266 452658 111502 452894
rect 111586 452658 111822 452894
rect 111266 452338 111502 452574
rect 111586 452338 111822 452574
rect 111266 418658 111502 418894
rect 111586 418658 111822 418894
rect 111266 418338 111502 418574
rect 111586 418338 111822 418574
rect 111266 384658 111502 384894
rect 111586 384658 111822 384894
rect 111266 384338 111502 384574
rect 111586 384338 111822 384574
rect 111266 350658 111502 350894
rect 111586 350658 111822 350894
rect 111266 350338 111502 350574
rect 111586 350338 111822 350574
rect 111266 316658 111502 316894
rect 111586 316658 111822 316894
rect 111266 316338 111502 316574
rect 111586 316338 111822 316574
rect 111266 282658 111502 282894
rect 111586 282658 111822 282894
rect 111266 282338 111502 282574
rect 111586 282338 111822 282574
rect 111266 248658 111502 248894
rect 111586 248658 111822 248894
rect 111266 248338 111502 248574
rect 111586 248338 111822 248574
rect 114986 707482 115222 707718
rect 115306 707482 115542 707718
rect 114986 707162 115222 707398
rect 115306 707162 115542 707398
rect 114986 694378 115222 694614
rect 115306 694378 115542 694614
rect 114986 694058 115222 694294
rect 115306 694058 115542 694294
rect 114986 660378 115222 660614
rect 115306 660378 115542 660614
rect 114986 660058 115222 660294
rect 115306 660058 115542 660294
rect 114986 626378 115222 626614
rect 115306 626378 115542 626614
rect 114986 626058 115222 626294
rect 115306 626058 115542 626294
rect 114986 592378 115222 592614
rect 115306 592378 115542 592614
rect 114986 592058 115222 592294
rect 115306 592058 115542 592294
rect 114986 558378 115222 558614
rect 115306 558378 115542 558614
rect 114986 558058 115222 558294
rect 115306 558058 115542 558294
rect 114986 524378 115222 524614
rect 115306 524378 115542 524614
rect 114986 524058 115222 524294
rect 115306 524058 115542 524294
rect 114986 490378 115222 490614
rect 115306 490378 115542 490614
rect 114986 490058 115222 490294
rect 115306 490058 115542 490294
rect 114986 456378 115222 456614
rect 115306 456378 115542 456614
rect 114986 456058 115222 456294
rect 115306 456058 115542 456294
rect 114986 422378 115222 422614
rect 115306 422378 115542 422614
rect 114986 422058 115222 422294
rect 115306 422058 115542 422294
rect 114986 388378 115222 388614
rect 115306 388378 115542 388614
rect 114986 388058 115222 388294
rect 115306 388058 115542 388294
rect 114986 354378 115222 354614
rect 115306 354378 115542 354614
rect 114986 354058 115222 354294
rect 115306 354058 115542 354294
rect 114986 320378 115222 320614
rect 115306 320378 115542 320614
rect 114986 320058 115222 320294
rect 115306 320058 115542 320294
rect 114986 286378 115222 286614
rect 115306 286378 115542 286614
rect 114986 286058 115222 286294
rect 115306 286058 115542 286294
rect 114986 252378 115222 252614
rect 115306 252378 115542 252614
rect 114986 252058 115222 252294
rect 115306 252058 115542 252294
rect 118706 708442 118942 708678
rect 119026 708442 119262 708678
rect 118706 708122 118942 708358
rect 119026 708122 119262 708358
rect 118706 698098 118942 698334
rect 119026 698098 119262 698334
rect 118706 697778 118942 698014
rect 119026 697778 119262 698014
rect 118706 664098 118942 664334
rect 119026 664098 119262 664334
rect 118706 663778 118942 664014
rect 119026 663778 119262 664014
rect 118706 630098 118942 630334
rect 119026 630098 119262 630334
rect 118706 629778 118942 630014
rect 119026 629778 119262 630014
rect 118706 596098 118942 596334
rect 119026 596098 119262 596334
rect 118706 595778 118942 596014
rect 119026 595778 119262 596014
rect 118706 562098 118942 562334
rect 119026 562098 119262 562334
rect 118706 561778 118942 562014
rect 119026 561778 119262 562014
rect 118706 528098 118942 528334
rect 119026 528098 119262 528334
rect 118706 527778 118942 528014
rect 119026 527778 119262 528014
rect 118706 494098 118942 494334
rect 119026 494098 119262 494334
rect 118706 493778 118942 494014
rect 119026 493778 119262 494014
rect 118706 460098 118942 460334
rect 119026 460098 119262 460334
rect 118706 459778 118942 460014
rect 119026 459778 119262 460014
rect 118706 426098 118942 426334
rect 119026 426098 119262 426334
rect 118706 425778 118942 426014
rect 119026 425778 119262 426014
rect 118706 392098 118942 392334
rect 119026 392098 119262 392334
rect 118706 391778 118942 392014
rect 119026 391778 119262 392014
rect 118706 358098 118942 358334
rect 119026 358098 119262 358334
rect 118706 357778 118942 358014
rect 119026 357778 119262 358014
rect 118706 324098 118942 324334
rect 119026 324098 119262 324334
rect 118706 323778 118942 324014
rect 119026 323778 119262 324014
rect 118706 290098 118942 290334
rect 119026 290098 119262 290334
rect 118706 289778 118942 290014
rect 119026 289778 119262 290014
rect 118706 256098 118942 256334
rect 119026 256098 119262 256334
rect 118706 255778 118942 256014
rect 119026 255778 119262 256014
rect 122426 709402 122662 709638
rect 122746 709402 122982 709638
rect 122426 709082 122662 709318
rect 122746 709082 122982 709318
rect 122426 667818 122662 668054
rect 122746 667818 122982 668054
rect 122426 667498 122662 667734
rect 122746 667498 122982 667734
rect 122426 633818 122662 634054
rect 122746 633818 122982 634054
rect 122426 633498 122662 633734
rect 122746 633498 122982 633734
rect 122426 599818 122662 600054
rect 122746 599818 122982 600054
rect 122426 599498 122662 599734
rect 122746 599498 122982 599734
rect 122426 565818 122662 566054
rect 122746 565818 122982 566054
rect 122426 565498 122662 565734
rect 122746 565498 122982 565734
rect 122426 531818 122662 532054
rect 122746 531818 122982 532054
rect 122426 531498 122662 531734
rect 122746 531498 122982 531734
rect 122426 497818 122662 498054
rect 122746 497818 122982 498054
rect 122426 497498 122662 497734
rect 122746 497498 122982 497734
rect 122426 463818 122662 464054
rect 122746 463818 122982 464054
rect 122426 463498 122662 463734
rect 122746 463498 122982 463734
rect 122426 429818 122662 430054
rect 122746 429818 122982 430054
rect 122426 429498 122662 429734
rect 122746 429498 122982 429734
rect 122426 395818 122662 396054
rect 122746 395818 122982 396054
rect 122426 395498 122662 395734
rect 122746 395498 122982 395734
rect 122426 361818 122662 362054
rect 122746 361818 122982 362054
rect 122426 361498 122662 361734
rect 122746 361498 122982 361734
rect 122426 327818 122662 328054
rect 122746 327818 122982 328054
rect 122426 327498 122662 327734
rect 122746 327498 122982 327734
rect 122426 293818 122662 294054
rect 122746 293818 122982 294054
rect 122426 293498 122662 293734
rect 122746 293498 122982 293734
rect 122426 259818 122662 260054
rect 122746 259818 122982 260054
rect 122426 259498 122662 259734
rect 122746 259498 122982 259734
rect 122426 225755 122662 225991
rect 122746 225755 122982 225991
rect 126146 710362 126382 710598
rect 126466 710362 126702 710598
rect 126146 710042 126382 710278
rect 126466 710042 126702 710278
rect 126146 671538 126382 671774
rect 126466 671538 126702 671774
rect 126146 671218 126382 671454
rect 126466 671218 126702 671454
rect 126146 637538 126382 637774
rect 126466 637538 126702 637774
rect 126146 637218 126382 637454
rect 126466 637218 126702 637454
rect 126146 603538 126382 603774
rect 126466 603538 126702 603774
rect 126146 603218 126382 603454
rect 126466 603218 126702 603454
rect 126146 569538 126382 569774
rect 126466 569538 126702 569774
rect 126146 569218 126382 569454
rect 126466 569218 126702 569454
rect 126146 535538 126382 535774
rect 126466 535538 126702 535774
rect 126146 535218 126382 535454
rect 126466 535218 126702 535454
rect 126146 501538 126382 501774
rect 126466 501538 126702 501774
rect 126146 501218 126382 501454
rect 126466 501218 126702 501454
rect 126146 467538 126382 467774
rect 126466 467538 126702 467774
rect 126146 467218 126382 467454
rect 126466 467218 126702 467454
rect 126146 433538 126382 433774
rect 126466 433538 126702 433774
rect 126146 433218 126382 433454
rect 126466 433218 126702 433454
rect 126146 399538 126382 399774
rect 126466 399538 126702 399774
rect 126146 399218 126382 399454
rect 126466 399218 126702 399454
rect 126146 365538 126382 365774
rect 126466 365538 126702 365774
rect 126146 365218 126382 365454
rect 126466 365218 126702 365454
rect 126146 331538 126382 331774
rect 126466 331538 126702 331774
rect 126146 331218 126382 331454
rect 126466 331218 126702 331454
rect 126146 297538 126382 297774
rect 126466 297538 126702 297774
rect 126146 297218 126382 297454
rect 126466 297218 126702 297454
rect 126146 263538 126382 263774
rect 126466 263538 126702 263774
rect 126146 263218 126382 263454
rect 126466 263218 126702 263454
rect 126146 229538 126382 229774
rect 126466 229538 126702 229774
rect 126146 229218 126382 229454
rect 126466 229218 126702 229454
rect 129866 711322 130102 711558
rect 130186 711322 130422 711558
rect 129866 711002 130102 711238
rect 130186 711002 130422 711238
rect 129866 675258 130102 675494
rect 130186 675258 130422 675494
rect 129866 674938 130102 675174
rect 130186 674938 130422 675174
rect 129866 641258 130102 641494
rect 130186 641258 130422 641494
rect 129866 640938 130102 641174
rect 130186 640938 130422 641174
rect 129866 607258 130102 607494
rect 130186 607258 130422 607494
rect 129866 606938 130102 607174
rect 130186 606938 130422 607174
rect 129866 573258 130102 573494
rect 130186 573258 130422 573494
rect 129866 572938 130102 573174
rect 130186 572938 130422 573174
rect 129866 539258 130102 539494
rect 130186 539258 130422 539494
rect 129866 538938 130102 539174
rect 130186 538938 130422 539174
rect 129866 505258 130102 505494
rect 130186 505258 130422 505494
rect 129866 504938 130102 505174
rect 130186 504938 130422 505174
rect 129866 471258 130102 471494
rect 130186 471258 130422 471494
rect 129866 470938 130102 471174
rect 130186 470938 130422 471174
rect 129866 437258 130102 437494
rect 130186 437258 130422 437494
rect 129866 436938 130102 437174
rect 130186 436938 130422 437174
rect 129866 403258 130102 403494
rect 130186 403258 130422 403494
rect 129866 402938 130102 403174
rect 130186 402938 130422 403174
rect 129866 369258 130102 369494
rect 130186 369258 130422 369494
rect 129866 368938 130102 369174
rect 130186 368938 130422 369174
rect 129866 335258 130102 335494
rect 130186 335258 130422 335494
rect 129866 334938 130102 335174
rect 130186 334938 130422 335174
rect 129866 301258 130102 301494
rect 130186 301258 130422 301494
rect 129866 300938 130102 301174
rect 130186 300938 130422 301174
rect 129866 267258 130102 267494
rect 130186 267258 130422 267494
rect 129866 266938 130102 267174
rect 130186 266938 130422 267174
rect 129866 233258 130102 233494
rect 130186 233258 130422 233494
rect 129866 232938 130102 233174
rect 130186 232938 130422 233174
rect 43266 214658 43502 214894
rect 43586 214658 43822 214894
rect 43266 214338 43502 214574
rect 43586 214338 43822 214574
rect 43266 180658 43502 180894
rect 43586 180658 43822 180894
rect 43266 180338 43502 180574
rect 43586 180338 43822 180574
rect 43266 146658 43502 146894
rect 43586 146658 43822 146894
rect 43266 146338 43502 146574
rect 43586 146338 43822 146574
rect 43266 112658 43502 112894
rect 43586 112658 43822 112894
rect 43266 112338 43502 112574
rect 43586 112338 43822 112574
rect 43266 78658 43502 78894
rect 43586 78658 43822 78894
rect 43266 78338 43502 78574
rect 43586 78338 43822 78574
rect 43266 44658 43502 44894
rect 43586 44658 43822 44894
rect 43266 44338 43502 44574
rect 43586 44338 43822 44574
rect 43266 10658 43502 10894
rect 43586 10658 43822 10894
rect 43266 10338 43502 10574
rect 43586 10338 43822 10574
rect 43266 -2502 43502 -2266
rect 43586 -2502 43822 -2266
rect 43266 -2822 43502 -2586
rect 43586 -2822 43822 -2586
rect 46986 184378 47222 184614
rect 47306 184378 47542 184614
rect 46986 184058 47222 184294
rect 47306 184058 47542 184294
rect 46986 150378 47222 150614
rect 47306 150378 47542 150614
rect 46986 150058 47222 150294
rect 47306 150058 47542 150294
rect 46986 116378 47222 116614
rect 47306 116378 47542 116614
rect 46986 116058 47222 116294
rect 47306 116058 47542 116294
rect 46986 82378 47222 82614
rect 47306 82378 47542 82614
rect 46986 82058 47222 82294
rect 47306 82058 47542 82294
rect 46986 48378 47222 48614
rect 47306 48378 47542 48614
rect 46986 48058 47222 48294
rect 47306 48058 47542 48294
rect 46986 14378 47222 14614
rect 47306 14378 47542 14614
rect 46986 14058 47222 14294
rect 47306 14058 47542 14294
rect 46986 -3462 47222 -3226
rect 47306 -3462 47542 -3226
rect 46986 -3782 47222 -3546
rect 47306 -3782 47542 -3546
rect 50706 188098 50942 188334
rect 51026 188098 51262 188334
rect 50706 187778 50942 188014
rect 51026 187778 51262 188014
rect 50706 154098 50942 154334
rect 51026 154098 51262 154334
rect 50706 153778 50942 154014
rect 51026 153778 51262 154014
rect 50706 120098 50942 120334
rect 51026 120098 51262 120334
rect 50706 119778 50942 120014
rect 51026 119778 51262 120014
rect 50706 86098 50942 86334
rect 51026 86098 51262 86334
rect 50706 85778 50942 86014
rect 51026 85778 51262 86014
rect 50706 52098 50942 52334
rect 51026 52098 51262 52334
rect 50706 51778 50942 52014
rect 51026 51778 51262 52014
rect 50706 18098 50942 18334
rect 51026 18098 51262 18334
rect 50706 17778 50942 18014
rect 51026 17778 51262 18014
rect 50706 -4422 50942 -4186
rect 51026 -4422 51262 -4186
rect 50706 -4742 50942 -4506
rect 51026 -4742 51262 -4506
rect 54426 191818 54662 192054
rect 54746 191818 54982 192054
rect 54426 191498 54662 191734
rect 54746 191498 54982 191734
rect 54426 157818 54662 158054
rect 54746 157818 54982 158054
rect 54426 157498 54662 157734
rect 54746 157498 54982 157734
rect 54426 123818 54662 124054
rect 54746 123818 54982 124054
rect 54426 123498 54662 123734
rect 54746 123498 54982 123734
rect 54426 89818 54662 90054
rect 54746 89818 54982 90054
rect 54426 89498 54662 89734
rect 54746 89498 54982 89734
rect 54426 55818 54662 56054
rect 54746 55818 54982 56054
rect 54426 55498 54662 55734
rect 54746 55498 54982 55734
rect 54426 21818 54662 22054
rect 54746 21818 54982 22054
rect 54426 21498 54662 21734
rect 54746 21498 54982 21734
rect 54426 -5382 54662 -5146
rect 54746 -5382 54982 -5146
rect 54426 -5702 54662 -5466
rect 54746 -5702 54982 -5466
rect 58146 195538 58382 195774
rect 58466 195538 58702 195774
rect 58146 195218 58382 195454
rect 58466 195218 58702 195454
rect 58146 161538 58382 161774
rect 58466 161538 58702 161774
rect 58146 161218 58382 161454
rect 58466 161218 58702 161454
rect 58146 127538 58382 127774
rect 58466 127538 58702 127774
rect 58146 127218 58382 127454
rect 58466 127218 58702 127454
rect 58146 93538 58382 93774
rect 58466 93538 58702 93774
rect 58146 93218 58382 93454
rect 58466 93218 58702 93454
rect 58146 59538 58382 59774
rect 58466 59538 58702 59774
rect 58146 59218 58382 59454
rect 58466 59218 58702 59454
rect 58146 25538 58382 25774
rect 58466 25538 58702 25774
rect 58146 25218 58382 25454
rect 58466 25218 58702 25454
rect 58146 -6342 58382 -6106
rect 58466 -6342 58702 -6106
rect 58146 -6662 58382 -6426
rect 58466 -6662 58702 -6426
rect 61866 199258 62102 199494
rect 62186 199258 62422 199494
rect 61866 198938 62102 199174
rect 62186 198938 62422 199174
rect 61866 165258 62102 165494
rect 62186 165258 62422 165494
rect 61866 164938 62102 165174
rect 62186 164938 62422 165174
rect 61866 131258 62102 131494
rect 62186 131258 62422 131494
rect 61866 130938 62102 131174
rect 62186 130938 62422 131174
rect 61866 97258 62102 97494
rect 62186 97258 62422 97494
rect 61866 96938 62102 97174
rect 62186 96938 62422 97174
rect 61866 63258 62102 63494
rect 62186 63258 62422 63494
rect 61866 62938 62102 63174
rect 62186 62938 62422 63174
rect 61866 29258 62102 29494
rect 62186 29258 62422 29494
rect 61866 28938 62102 29174
rect 62186 28938 62422 29174
rect 61866 -7302 62102 -7066
rect 62186 -7302 62422 -7066
rect 61866 -7622 62102 -7386
rect 62186 -7622 62422 -7386
rect 69826 207218 70062 207454
rect 70146 207218 70382 207454
rect 69826 206898 70062 207134
rect 70146 206898 70382 207134
rect 69826 173218 70062 173454
rect 70146 173218 70382 173454
rect 69826 172898 70062 173134
rect 70146 172898 70382 173134
rect 69826 139218 70062 139454
rect 70146 139218 70382 139454
rect 69826 138898 70062 139134
rect 70146 138898 70382 139134
rect 69826 105218 70062 105454
rect 70146 105218 70382 105454
rect 69826 104898 70062 105134
rect 70146 104898 70382 105134
rect 69826 71218 70062 71454
rect 70146 71218 70382 71454
rect 69826 70898 70062 71134
rect 70146 70898 70382 71134
rect 69826 37218 70062 37454
rect 70146 37218 70382 37454
rect 69826 36898 70062 37134
rect 70146 36898 70382 37134
rect 69826 3218 70062 3454
rect 70146 3218 70382 3454
rect 69826 2898 70062 3134
rect 70146 2898 70382 3134
rect 69826 -582 70062 -346
rect 70146 -582 70382 -346
rect 69826 -902 70062 -666
rect 70146 -902 70382 -666
rect 73546 210938 73782 211174
rect 73866 210938 74102 211174
rect 73546 210618 73782 210854
rect 73866 210618 74102 210854
rect 73546 176938 73782 177174
rect 73866 176938 74102 177174
rect 73546 176618 73782 176854
rect 73866 176618 74102 176854
rect 73546 142938 73782 143174
rect 73866 142938 74102 143174
rect 73546 142618 73782 142854
rect 73866 142618 74102 142854
rect 73546 108938 73782 109174
rect 73866 108938 74102 109174
rect 73546 108618 73782 108854
rect 73866 108618 74102 108854
rect 73546 74938 73782 75174
rect 73866 74938 74102 75174
rect 73546 74618 73782 74854
rect 73866 74618 74102 74854
rect 73546 40938 73782 41174
rect 73866 40938 74102 41174
rect 73546 40618 73782 40854
rect 73866 40618 74102 40854
rect 73546 6938 73782 7174
rect 73866 6938 74102 7174
rect 73546 6618 73782 6854
rect 73866 6618 74102 6854
rect 73546 -1542 73782 -1306
rect 73866 -1542 74102 -1306
rect 73546 -1862 73782 -1626
rect 73866 -1862 74102 -1626
rect 77266 180658 77502 180894
rect 77586 180658 77822 180894
rect 77266 180338 77502 180574
rect 77586 180338 77822 180574
rect 77266 146658 77502 146894
rect 77586 146658 77822 146894
rect 77266 146338 77502 146574
rect 77586 146338 77822 146574
rect 77266 112658 77502 112894
rect 77586 112658 77822 112894
rect 77266 112338 77502 112574
rect 77586 112338 77822 112574
rect 77266 78658 77502 78894
rect 77586 78658 77822 78894
rect 77266 78338 77502 78574
rect 77586 78338 77822 78574
rect 77266 44658 77502 44894
rect 77586 44658 77822 44894
rect 77266 44338 77502 44574
rect 77586 44338 77822 44574
rect 77266 10658 77502 10894
rect 77586 10658 77822 10894
rect 77266 10338 77502 10574
rect 77586 10338 77822 10574
rect 77266 -2502 77502 -2266
rect 77586 -2502 77822 -2266
rect 77266 -2822 77502 -2586
rect 77586 -2822 77822 -2586
rect 80986 184378 81222 184614
rect 81306 184378 81542 184614
rect 80986 184058 81222 184294
rect 81306 184058 81542 184294
rect 80986 150378 81222 150614
rect 81306 150378 81542 150614
rect 80986 150058 81222 150294
rect 81306 150058 81542 150294
rect 80986 116378 81222 116614
rect 81306 116378 81542 116614
rect 80986 116058 81222 116294
rect 81306 116058 81542 116294
rect 80986 82378 81222 82614
rect 81306 82378 81542 82614
rect 80986 82058 81222 82294
rect 81306 82058 81542 82294
rect 80986 48378 81222 48614
rect 81306 48378 81542 48614
rect 80986 48058 81222 48294
rect 81306 48058 81542 48294
rect 80986 14378 81222 14614
rect 81306 14378 81542 14614
rect 80986 14058 81222 14294
rect 81306 14058 81542 14294
rect 80986 -3462 81222 -3226
rect 81306 -3462 81542 -3226
rect 80986 -3782 81222 -3546
rect 81306 -3782 81542 -3546
rect 84706 188098 84942 188334
rect 85026 188098 85262 188334
rect 84706 187778 84942 188014
rect 85026 187778 85262 188014
rect 84706 154098 84942 154334
rect 85026 154098 85262 154334
rect 84706 153778 84942 154014
rect 85026 153778 85262 154014
rect 84706 120098 84942 120334
rect 85026 120098 85262 120334
rect 84706 119778 84942 120014
rect 85026 119778 85262 120014
rect 84706 86098 84942 86334
rect 85026 86098 85262 86334
rect 84706 85778 84942 86014
rect 85026 85778 85262 86014
rect 84706 52098 84942 52334
rect 85026 52098 85262 52334
rect 84706 51778 84942 52014
rect 85026 51778 85262 52014
rect 84706 18098 84942 18334
rect 85026 18098 85262 18334
rect 84706 17778 84942 18014
rect 85026 17778 85262 18014
rect 84706 -4422 84942 -4186
rect 85026 -4422 85262 -4186
rect 84706 -4742 84942 -4506
rect 85026 -4742 85262 -4506
rect 88426 191818 88662 192054
rect 88746 191818 88982 192054
rect 88426 191498 88662 191734
rect 88746 191498 88982 191734
rect 88426 157818 88662 158054
rect 88746 157818 88982 158054
rect 88426 157498 88662 157734
rect 88746 157498 88982 157734
rect 88426 123818 88662 124054
rect 88746 123818 88982 124054
rect 88426 123498 88662 123734
rect 88746 123498 88982 123734
rect 88426 89818 88662 90054
rect 88746 89818 88982 90054
rect 88426 89498 88662 89734
rect 88746 89498 88982 89734
rect 88426 55818 88662 56054
rect 88746 55818 88982 56054
rect 88426 55498 88662 55734
rect 88746 55498 88982 55734
rect 88426 21818 88662 22054
rect 88746 21818 88982 22054
rect 88426 21498 88662 21734
rect 88746 21498 88982 21734
rect 88426 -5382 88662 -5146
rect 88746 -5382 88982 -5146
rect 88426 -5702 88662 -5466
rect 88746 -5702 88982 -5466
rect 92146 195538 92382 195774
rect 92466 195538 92702 195774
rect 92146 195218 92382 195454
rect 92466 195218 92702 195454
rect 92146 161538 92382 161774
rect 92466 161538 92702 161774
rect 92146 161218 92382 161454
rect 92466 161218 92702 161454
rect 92146 127538 92382 127774
rect 92466 127538 92702 127774
rect 92146 127218 92382 127454
rect 92466 127218 92702 127454
rect 92146 93538 92382 93774
rect 92466 93538 92702 93774
rect 92146 93218 92382 93454
rect 92466 93218 92702 93454
rect 92146 59538 92382 59774
rect 92466 59538 92702 59774
rect 92146 59218 92382 59454
rect 92466 59218 92702 59454
rect 92146 25538 92382 25774
rect 92466 25538 92702 25774
rect 92146 25218 92382 25454
rect 92466 25218 92702 25454
rect 92146 -6342 92382 -6106
rect 92466 -6342 92702 -6106
rect 92146 -6662 92382 -6426
rect 92466 -6662 92702 -6426
rect 95866 199258 96102 199494
rect 96186 199258 96422 199494
rect 95866 198938 96102 199174
rect 96186 198938 96422 199174
rect 95866 165258 96102 165494
rect 96186 165258 96422 165494
rect 95866 164938 96102 165174
rect 96186 164938 96422 165174
rect 95866 131258 96102 131494
rect 96186 131258 96422 131494
rect 95866 130938 96102 131174
rect 96186 130938 96422 131174
rect 95866 97258 96102 97494
rect 96186 97258 96422 97494
rect 95866 96938 96102 97174
rect 96186 96938 96422 97174
rect 95866 63258 96102 63494
rect 96186 63258 96422 63494
rect 95866 62938 96102 63174
rect 96186 62938 96422 63174
rect 95866 29258 96102 29494
rect 96186 29258 96422 29494
rect 95866 28938 96102 29174
rect 96186 28938 96422 29174
rect 95866 -7302 96102 -7066
rect 96186 -7302 96422 -7066
rect 95866 -7622 96102 -7386
rect 96186 -7622 96422 -7386
rect 103826 207218 104062 207454
rect 104146 207218 104382 207454
rect 103826 206898 104062 207134
rect 104146 206898 104382 207134
rect 103826 173218 104062 173454
rect 104146 173218 104382 173454
rect 103826 172898 104062 173134
rect 104146 172898 104382 173134
rect 103826 139218 104062 139454
rect 104146 139218 104382 139454
rect 103826 138898 104062 139134
rect 104146 138898 104382 139134
rect 103826 105218 104062 105454
rect 104146 105218 104382 105454
rect 103826 104898 104062 105134
rect 104146 104898 104382 105134
rect 103826 71218 104062 71454
rect 104146 71218 104382 71454
rect 103826 70898 104062 71134
rect 104146 70898 104382 71134
rect 103826 37218 104062 37454
rect 104146 37218 104382 37454
rect 103826 36898 104062 37134
rect 104146 36898 104382 37134
rect 103826 3218 104062 3454
rect 104146 3218 104382 3454
rect 103826 2898 104062 3134
rect 104146 2898 104382 3134
rect 103826 -582 104062 -346
rect 104146 -582 104382 -346
rect 103826 -902 104062 -666
rect 104146 -902 104382 -666
rect 107546 210938 107782 211174
rect 107866 210938 108102 211174
rect 107546 210618 107782 210854
rect 107866 210618 108102 210854
rect 107546 176938 107782 177174
rect 107866 176938 108102 177174
rect 107546 176618 107782 176854
rect 107866 176618 108102 176854
rect 107546 142938 107782 143174
rect 107866 142938 108102 143174
rect 107546 142618 107782 142854
rect 107866 142618 108102 142854
rect 107546 108938 107782 109174
rect 107866 108938 108102 109174
rect 107546 108618 107782 108854
rect 107866 108618 108102 108854
rect 107546 74938 107782 75174
rect 107866 74938 108102 75174
rect 107546 74618 107782 74854
rect 107866 74618 108102 74854
rect 107546 40938 107782 41174
rect 107866 40938 108102 41174
rect 107546 40618 107782 40854
rect 107866 40618 108102 40854
rect 107546 6938 107782 7174
rect 107866 6938 108102 7174
rect 107546 6618 107782 6854
rect 107866 6618 108102 6854
rect 107546 -1542 107782 -1306
rect 107866 -1542 108102 -1306
rect 107546 -1862 107782 -1626
rect 107866 -1862 108102 -1626
rect 111266 180658 111502 180894
rect 111586 180658 111822 180894
rect 111266 180338 111502 180574
rect 111586 180338 111822 180574
rect 111266 146658 111502 146894
rect 111586 146658 111822 146894
rect 111266 146338 111502 146574
rect 111586 146338 111822 146574
rect 111266 112658 111502 112894
rect 111586 112658 111822 112894
rect 111266 112338 111502 112574
rect 111586 112338 111822 112574
rect 111266 78658 111502 78894
rect 111586 78658 111822 78894
rect 111266 78338 111502 78574
rect 111586 78338 111822 78574
rect 111266 44658 111502 44894
rect 111586 44658 111822 44894
rect 111266 44338 111502 44574
rect 111586 44338 111822 44574
rect 111266 10658 111502 10894
rect 111586 10658 111822 10894
rect 111266 10338 111502 10574
rect 111586 10338 111822 10574
rect 111266 -2502 111502 -2266
rect 111586 -2502 111822 -2266
rect 111266 -2822 111502 -2586
rect 111586 -2822 111822 -2586
rect 114986 184378 115222 184614
rect 115306 184378 115542 184614
rect 114986 184058 115222 184294
rect 115306 184058 115542 184294
rect 114986 150378 115222 150614
rect 115306 150378 115542 150614
rect 114986 150058 115222 150294
rect 115306 150058 115542 150294
rect 118706 188098 118942 188334
rect 119026 188098 119262 188334
rect 118706 187778 118942 188014
rect 119026 187778 119262 188014
rect 118706 154098 118942 154334
rect 119026 154098 119262 154334
rect 118706 153778 118942 154014
rect 119026 153778 119262 154014
rect 122426 191818 122662 192054
rect 122746 191818 122982 192054
rect 122426 191498 122662 191734
rect 122746 191498 122982 191734
rect 122426 157818 122662 158054
rect 122746 157818 122982 158054
rect 122426 157498 122662 157734
rect 122746 157498 122982 157734
rect 126146 195538 126382 195774
rect 126466 195538 126702 195774
rect 126146 195218 126382 195454
rect 126466 195218 126702 195454
rect 126146 161538 126382 161774
rect 126466 161538 126702 161774
rect 126146 161218 126382 161454
rect 126466 161218 126702 161454
rect 137826 704602 138062 704838
rect 138146 704602 138382 704838
rect 137826 704282 138062 704518
rect 138146 704282 138382 704518
rect 137826 683218 138062 683454
rect 138146 683218 138382 683454
rect 137826 682898 138062 683134
rect 138146 682898 138382 683134
rect 137826 649218 138062 649454
rect 138146 649218 138382 649454
rect 137826 648898 138062 649134
rect 138146 648898 138382 649134
rect 137826 615218 138062 615454
rect 138146 615218 138382 615454
rect 137826 614898 138062 615134
rect 138146 614898 138382 615134
rect 137826 581218 138062 581454
rect 138146 581218 138382 581454
rect 137826 580898 138062 581134
rect 138146 580898 138382 581134
rect 137826 547218 138062 547454
rect 138146 547218 138382 547454
rect 137826 546898 138062 547134
rect 138146 546898 138382 547134
rect 137826 513218 138062 513454
rect 138146 513218 138382 513454
rect 137826 512898 138062 513134
rect 138146 512898 138382 513134
rect 137826 479218 138062 479454
rect 138146 479218 138382 479454
rect 137826 478898 138062 479134
rect 138146 478898 138382 479134
rect 137826 445218 138062 445454
rect 138146 445218 138382 445454
rect 137826 444898 138062 445134
rect 138146 444898 138382 445134
rect 137826 411218 138062 411454
rect 138146 411218 138382 411454
rect 137826 410898 138062 411134
rect 138146 410898 138382 411134
rect 137826 377218 138062 377454
rect 138146 377218 138382 377454
rect 137826 376898 138062 377134
rect 138146 376898 138382 377134
rect 137826 343218 138062 343454
rect 138146 343218 138382 343454
rect 137826 342898 138062 343134
rect 138146 342898 138382 343134
rect 137826 309218 138062 309454
rect 138146 309218 138382 309454
rect 137826 308898 138062 309134
rect 138146 308898 138382 309134
rect 137826 275218 138062 275454
rect 138146 275218 138382 275454
rect 137826 274898 138062 275134
rect 138146 274898 138382 275134
rect 137826 241218 138062 241454
rect 138146 241218 138382 241454
rect 137826 240898 138062 241134
rect 138146 240898 138382 241134
rect 141546 705562 141782 705798
rect 141866 705562 142102 705798
rect 141546 705242 141782 705478
rect 141866 705242 142102 705478
rect 141546 686938 141782 687174
rect 141866 686938 142102 687174
rect 141546 686618 141782 686854
rect 141866 686618 142102 686854
rect 141546 652938 141782 653174
rect 141866 652938 142102 653174
rect 141546 652618 141782 652854
rect 141866 652618 142102 652854
rect 141546 618938 141782 619174
rect 141866 618938 142102 619174
rect 141546 618618 141782 618854
rect 141866 618618 142102 618854
rect 141546 584938 141782 585174
rect 141866 584938 142102 585174
rect 141546 584618 141782 584854
rect 141866 584618 142102 584854
rect 141546 550938 141782 551174
rect 141866 550938 142102 551174
rect 141546 550618 141782 550854
rect 141866 550618 142102 550854
rect 141546 516938 141782 517174
rect 141866 516938 142102 517174
rect 141546 516618 141782 516854
rect 141866 516618 142102 516854
rect 141546 482938 141782 483174
rect 141866 482938 142102 483174
rect 141546 482618 141782 482854
rect 141866 482618 142102 482854
rect 141546 448938 141782 449174
rect 141866 448938 142102 449174
rect 141546 448618 141782 448854
rect 141866 448618 142102 448854
rect 141546 414938 141782 415174
rect 141866 414938 142102 415174
rect 141546 414618 141782 414854
rect 141866 414618 142102 414854
rect 141546 380938 141782 381174
rect 141866 380938 142102 381174
rect 141546 380618 141782 380854
rect 141866 380618 142102 380854
rect 141546 346938 141782 347174
rect 141866 346938 142102 347174
rect 141546 346618 141782 346854
rect 141866 346618 142102 346854
rect 141546 312938 141782 313174
rect 141866 312938 142102 313174
rect 141546 312618 141782 312854
rect 141866 312618 142102 312854
rect 141546 278938 141782 279174
rect 141866 278938 142102 279174
rect 141546 278618 141782 278854
rect 141866 278618 142102 278854
rect 141546 244938 141782 245174
rect 141866 244938 142102 245174
rect 141546 244618 141782 244854
rect 141866 244618 142102 244854
rect 145266 706522 145502 706758
rect 145586 706522 145822 706758
rect 145266 706202 145502 706438
rect 145586 706202 145822 706438
rect 145266 690658 145502 690894
rect 145586 690658 145822 690894
rect 145266 690338 145502 690574
rect 145586 690338 145822 690574
rect 145266 656658 145502 656894
rect 145586 656658 145822 656894
rect 145266 656338 145502 656574
rect 145586 656338 145822 656574
rect 145266 622658 145502 622894
rect 145586 622658 145822 622894
rect 145266 622338 145502 622574
rect 145586 622338 145822 622574
rect 145266 588658 145502 588894
rect 145586 588658 145822 588894
rect 145266 588338 145502 588574
rect 145586 588338 145822 588574
rect 145266 554658 145502 554894
rect 145586 554658 145822 554894
rect 145266 554338 145502 554574
rect 145586 554338 145822 554574
rect 145266 520658 145502 520894
rect 145586 520658 145822 520894
rect 145266 520338 145502 520574
rect 145586 520338 145822 520574
rect 145266 486658 145502 486894
rect 145586 486658 145822 486894
rect 145266 486338 145502 486574
rect 145586 486338 145822 486574
rect 145266 452658 145502 452894
rect 145586 452658 145822 452894
rect 145266 452338 145502 452574
rect 145586 452338 145822 452574
rect 145266 418658 145502 418894
rect 145586 418658 145822 418894
rect 145266 418338 145502 418574
rect 145586 418338 145822 418574
rect 145266 384658 145502 384894
rect 145586 384658 145822 384894
rect 145266 384338 145502 384574
rect 145586 384338 145822 384574
rect 145266 350658 145502 350894
rect 145586 350658 145822 350894
rect 145266 350338 145502 350574
rect 145586 350338 145822 350574
rect 145266 316658 145502 316894
rect 145586 316658 145822 316894
rect 145266 316338 145502 316574
rect 145586 316338 145822 316574
rect 145266 282658 145502 282894
rect 145586 282658 145822 282894
rect 145266 282338 145502 282574
rect 145586 282338 145822 282574
rect 145266 248658 145502 248894
rect 145586 248658 145822 248894
rect 145266 248338 145502 248574
rect 145586 248338 145822 248574
rect 148986 707482 149222 707718
rect 149306 707482 149542 707718
rect 148986 707162 149222 707398
rect 149306 707162 149542 707398
rect 148986 694378 149222 694614
rect 149306 694378 149542 694614
rect 148986 694058 149222 694294
rect 149306 694058 149542 694294
rect 148986 660378 149222 660614
rect 149306 660378 149542 660614
rect 148986 660058 149222 660294
rect 149306 660058 149542 660294
rect 148986 626378 149222 626614
rect 149306 626378 149542 626614
rect 148986 626058 149222 626294
rect 149306 626058 149542 626294
rect 148986 592378 149222 592614
rect 149306 592378 149542 592614
rect 148986 592058 149222 592294
rect 149306 592058 149542 592294
rect 148986 558378 149222 558614
rect 149306 558378 149542 558614
rect 148986 558058 149222 558294
rect 149306 558058 149542 558294
rect 148986 524378 149222 524614
rect 149306 524378 149542 524614
rect 148986 524058 149222 524294
rect 149306 524058 149542 524294
rect 148986 490378 149222 490614
rect 149306 490378 149542 490614
rect 148986 490058 149222 490294
rect 149306 490058 149542 490294
rect 148986 456378 149222 456614
rect 149306 456378 149542 456614
rect 148986 456058 149222 456294
rect 149306 456058 149542 456294
rect 148986 422378 149222 422614
rect 149306 422378 149542 422614
rect 148986 422058 149222 422294
rect 149306 422058 149542 422294
rect 148986 388378 149222 388614
rect 149306 388378 149542 388614
rect 148986 388058 149222 388294
rect 149306 388058 149542 388294
rect 148986 354378 149222 354614
rect 149306 354378 149542 354614
rect 148986 354058 149222 354294
rect 149306 354058 149542 354294
rect 148986 320378 149222 320614
rect 149306 320378 149542 320614
rect 148986 320058 149222 320294
rect 149306 320058 149542 320294
rect 148986 286378 149222 286614
rect 149306 286378 149542 286614
rect 148986 286058 149222 286294
rect 149306 286058 149542 286294
rect 148986 252378 149222 252614
rect 149306 252378 149542 252614
rect 148986 252058 149222 252294
rect 149306 252058 149542 252294
rect 152706 708442 152942 708678
rect 153026 708442 153262 708678
rect 152706 708122 152942 708358
rect 153026 708122 153262 708358
rect 152706 698098 152942 698334
rect 153026 698098 153262 698334
rect 152706 697778 152942 698014
rect 153026 697778 153262 698014
rect 152706 664098 152942 664334
rect 153026 664098 153262 664334
rect 152706 663778 152942 664014
rect 153026 663778 153262 664014
rect 152706 630098 152942 630334
rect 153026 630098 153262 630334
rect 152706 629778 152942 630014
rect 153026 629778 153262 630014
rect 152706 596098 152942 596334
rect 153026 596098 153262 596334
rect 152706 595778 152942 596014
rect 153026 595778 153262 596014
rect 152706 562098 152942 562334
rect 153026 562098 153262 562334
rect 152706 561778 152942 562014
rect 153026 561778 153262 562014
rect 152706 528098 152942 528334
rect 153026 528098 153262 528334
rect 152706 527778 152942 528014
rect 153026 527778 153262 528014
rect 152706 494098 152942 494334
rect 153026 494098 153262 494334
rect 152706 493778 152942 494014
rect 153026 493778 153262 494014
rect 152706 460098 152942 460334
rect 153026 460098 153262 460334
rect 152706 459778 152942 460014
rect 153026 459778 153262 460014
rect 152706 426098 152942 426334
rect 153026 426098 153262 426334
rect 152706 425778 152942 426014
rect 153026 425778 153262 426014
rect 152706 392098 152942 392334
rect 153026 392098 153262 392334
rect 152706 391778 152942 392014
rect 153026 391778 153262 392014
rect 152706 358098 152942 358334
rect 153026 358098 153262 358334
rect 152706 357778 152942 358014
rect 153026 357778 153262 358014
rect 152706 324098 152942 324334
rect 153026 324098 153262 324334
rect 152706 323778 152942 324014
rect 153026 323778 153262 324014
rect 152706 290098 152942 290334
rect 153026 290098 153262 290334
rect 152706 289778 152942 290014
rect 153026 289778 153262 290014
rect 152706 256098 152942 256334
rect 153026 256098 153262 256334
rect 152706 255778 152942 256014
rect 153026 255778 153262 256014
rect 156426 709402 156662 709638
rect 156746 709402 156982 709638
rect 156426 709082 156662 709318
rect 156746 709082 156982 709318
rect 156426 667818 156662 668054
rect 156746 667818 156982 668054
rect 156426 667498 156662 667734
rect 156746 667498 156982 667734
rect 156426 633818 156662 634054
rect 156746 633818 156982 634054
rect 156426 633498 156662 633734
rect 156746 633498 156982 633734
rect 156426 599818 156662 600054
rect 156746 599818 156982 600054
rect 156426 599498 156662 599734
rect 156746 599498 156982 599734
rect 156426 565818 156662 566054
rect 156746 565818 156982 566054
rect 156426 565498 156662 565734
rect 156746 565498 156982 565734
rect 156426 531818 156662 532054
rect 156746 531818 156982 532054
rect 156426 531498 156662 531734
rect 156746 531498 156982 531734
rect 156426 497818 156662 498054
rect 156746 497818 156982 498054
rect 156426 497498 156662 497734
rect 156746 497498 156982 497734
rect 156426 463818 156662 464054
rect 156746 463818 156982 464054
rect 156426 463498 156662 463734
rect 156746 463498 156982 463734
rect 156426 429818 156662 430054
rect 156746 429818 156982 430054
rect 156426 429498 156662 429734
rect 156746 429498 156982 429734
rect 156426 395818 156662 396054
rect 156746 395818 156982 396054
rect 156426 395498 156662 395734
rect 156746 395498 156982 395734
rect 156426 361818 156662 362054
rect 156746 361818 156982 362054
rect 156426 361498 156662 361734
rect 156746 361498 156982 361734
rect 156426 327818 156662 328054
rect 156746 327818 156982 328054
rect 156426 327498 156662 327734
rect 156746 327498 156982 327734
rect 156426 293818 156662 294054
rect 156746 293818 156982 294054
rect 156426 293498 156662 293734
rect 156746 293498 156982 293734
rect 156426 259818 156662 260054
rect 156746 259818 156982 260054
rect 156426 259498 156662 259734
rect 156746 259498 156982 259734
rect 156426 225755 156662 225991
rect 156746 225755 156982 225991
rect 160146 710362 160382 710598
rect 160466 710362 160702 710598
rect 160146 710042 160382 710278
rect 160466 710042 160702 710278
rect 160146 671538 160382 671774
rect 160466 671538 160702 671774
rect 160146 671218 160382 671454
rect 160466 671218 160702 671454
rect 160146 637538 160382 637774
rect 160466 637538 160702 637774
rect 160146 637218 160382 637454
rect 160466 637218 160702 637454
rect 160146 603538 160382 603774
rect 160466 603538 160702 603774
rect 160146 603218 160382 603454
rect 160466 603218 160702 603454
rect 160146 569538 160382 569774
rect 160466 569538 160702 569774
rect 160146 569218 160382 569454
rect 160466 569218 160702 569454
rect 160146 535538 160382 535774
rect 160466 535538 160702 535774
rect 160146 535218 160382 535454
rect 160466 535218 160702 535454
rect 160146 501538 160382 501774
rect 160466 501538 160702 501774
rect 160146 501218 160382 501454
rect 160466 501218 160702 501454
rect 160146 467538 160382 467774
rect 160466 467538 160702 467774
rect 160146 467218 160382 467454
rect 160466 467218 160702 467454
rect 160146 433538 160382 433774
rect 160466 433538 160702 433774
rect 160146 433218 160382 433454
rect 160466 433218 160702 433454
rect 160146 399538 160382 399774
rect 160466 399538 160702 399774
rect 160146 399218 160382 399454
rect 160466 399218 160702 399454
rect 160146 365538 160382 365774
rect 160466 365538 160702 365774
rect 160146 365218 160382 365454
rect 160466 365218 160702 365454
rect 160146 331538 160382 331774
rect 160466 331538 160702 331774
rect 160146 331218 160382 331454
rect 160466 331218 160702 331454
rect 160146 297538 160382 297774
rect 160466 297538 160702 297774
rect 160146 297218 160382 297454
rect 160466 297218 160702 297454
rect 160146 263538 160382 263774
rect 160466 263538 160702 263774
rect 160146 263218 160382 263454
rect 160466 263218 160702 263454
rect 160146 229538 160382 229774
rect 160466 229538 160702 229774
rect 160146 229218 160382 229454
rect 160466 229218 160702 229454
rect 129866 199258 130102 199494
rect 130186 199258 130422 199494
rect 129866 198938 130102 199174
rect 130186 198938 130422 199174
rect 163866 711322 164102 711558
rect 164186 711322 164422 711558
rect 163866 711002 164102 711238
rect 164186 711002 164422 711238
rect 163866 675258 164102 675494
rect 164186 675258 164422 675494
rect 163866 674938 164102 675174
rect 164186 674938 164422 675174
rect 163866 641258 164102 641494
rect 164186 641258 164422 641494
rect 163866 640938 164102 641174
rect 164186 640938 164422 641174
rect 163866 607258 164102 607494
rect 164186 607258 164422 607494
rect 163866 606938 164102 607174
rect 164186 606938 164422 607174
rect 163866 573258 164102 573494
rect 164186 573258 164422 573494
rect 163866 572938 164102 573174
rect 164186 572938 164422 573174
rect 163866 539258 164102 539494
rect 164186 539258 164422 539494
rect 163866 538938 164102 539174
rect 164186 538938 164422 539174
rect 163866 505258 164102 505494
rect 164186 505258 164422 505494
rect 163866 504938 164102 505174
rect 164186 504938 164422 505174
rect 163866 471258 164102 471494
rect 164186 471258 164422 471494
rect 163866 470938 164102 471174
rect 164186 470938 164422 471174
rect 163866 437258 164102 437494
rect 164186 437258 164422 437494
rect 163866 436938 164102 437174
rect 164186 436938 164422 437174
rect 163866 403258 164102 403494
rect 164186 403258 164422 403494
rect 163866 402938 164102 403174
rect 164186 402938 164422 403174
rect 163866 369258 164102 369494
rect 164186 369258 164422 369494
rect 163866 368938 164102 369174
rect 164186 368938 164422 369174
rect 163866 335258 164102 335494
rect 164186 335258 164422 335494
rect 163866 334938 164102 335174
rect 164186 334938 164422 335174
rect 163866 301258 164102 301494
rect 164186 301258 164422 301494
rect 163866 300938 164102 301174
rect 164186 300938 164422 301174
rect 163866 267258 164102 267494
rect 164186 267258 164422 267494
rect 163866 266938 164102 267174
rect 164186 266938 164422 267174
rect 163866 233258 164102 233494
rect 164186 233258 164422 233494
rect 163866 232938 164102 233174
rect 164186 232938 164422 233174
rect 171826 704602 172062 704838
rect 172146 704602 172382 704838
rect 171826 704282 172062 704518
rect 172146 704282 172382 704518
rect 171826 683218 172062 683454
rect 172146 683218 172382 683454
rect 171826 682898 172062 683134
rect 172146 682898 172382 683134
rect 171826 649218 172062 649454
rect 172146 649218 172382 649454
rect 171826 648898 172062 649134
rect 172146 648898 172382 649134
rect 171826 615218 172062 615454
rect 172146 615218 172382 615454
rect 171826 614898 172062 615134
rect 172146 614898 172382 615134
rect 171826 581218 172062 581454
rect 172146 581218 172382 581454
rect 171826 580898 172062 581134
rect 172146 580898 172382 581134
rect 171826 547218 172062 547454
rect 172146 547218 172382 547454
rect 171826 546898 172062 547134
rect 172146 546898 172382 547134
rect 171826 513218 172062 513454
rect 172146 513218 172382 513454
rect 171826 512898 172062 513134
rect 172146 512898 172382 513134
rect 171826 479218 172062 479454
rect 172146 479218 172382 479454
rect 171826 478898 172062 479134
rect 172146 478898 172382 479134
rect 171826 445218 172062 445454
rect 172146 445218 172382 445454
rect 171826 444898 172062 445134
rect 172146 444898 172382 445134
rect 171826 411218 172062 411454
rect 172146 411218 172382 411454
rect 171826 410898 172062 411134
rect 172146 410898 172382 411134
rect 171826 377218 172062 377454
rect 172146 377218 172382 377454
rect 171826 376898 172062 377134
rect 172146 376898 172382 377134
rect 171826 343218 172062 343454
rect 172146 343218 172382 343454
rect 171826 342898 172062 343134
rect 172146 342898 172382 343134
rect 171826 309218 172062 309454
rect 172146 309218 172382 309454
rect 171826 308898 172062 309134
rect 172146 308898 172382 309134
rect 171826 275218 172062 275454
rect 172146 275218 172382 275454
rect 171826 274898 172062 275134
rect 172146 274898 172382 275134
rect 171826 241218 172062 241454
rect 172146 241218 172382 241454
rect 171826 240898 172062 241134
rect 172146 240898 172382 241134
rect 175546 705562 175782 705798
rect 175866 705562 176102 705798
rect 175546 705242 175782 705478
rect 175866 705242 176102 705478
rect 175546 686938 175782 687174
rect 175866 686938 176102 687174
rect 175546 686618 175782 686854
rect 175866 686618 176102 686854
rect 175546 652938 175782 653174
rect 175866 652938 176102 653174
rect 175546 652618 175782 652854
rect 175866 652618 176102 652854
rect 175546 618938 175782 619174
rect 175866 618938 176102 619174
rect 175546 618618 175782 618854
rect 175866 618618 176102 618854
rect 175546 584938 175782 585174
rect 175866 584938 176102 585174
rect 175546 584618 175782 584854
rect 175866 584618 176102 584854
rect 175546 550938 175782 551174
rect 175866 550938 176102 551174
rect 175546 550618 175782 550854
rect 175866 550618 176102 550854
rect 175546 516938 175782 517174
rect 175866 516938 176102 517174
rect 175546 516618 175782 516854
rect 175866 516618 176102 516854
rect 175546 482938 175782 483174
rect 175866 482938 176102 483174
rect 175546 482618 175782 482854
rect 175866 482618 176102 482854
rect 175546 448938 175782 449174
rect 175866 448938 176102 449174
rect 175546 448618 175782 448854
rect 175866 448618 176102 448854
rect 175546 414938 175782 415174
rect 175866 414938 176102 415174
rect 175546 414618 175782 414854
rect 175866 414618 176102 414854
rect 175546 380938 175782 381174
rect 175866 380938 176102 381174
rect 175546 380618 175782 380854
rect 175866 380618 176102 380854
rect 175546 346938 175782 347174
rect 175866 346938 176102 347174
rect 175546 346618 175782 346854
rect 175866 346618 176102 346854
rect 175546 312938 175782 313174
rect 175866 312938 176102 313174
rect 175546 312618 175782 312854
rect 175866 312618 176102 312854
rect 175546 278938 175782 279174
rect 175866 278938 176102 279174
rect 175546 278618 175782 278854
rect 175866 278618 176102 278854
rect 175546 244938 175782 245174
rect 175866 244938 176102 245174
rect 175546 244618 175782 244854
rect 175866 244618 176102 244854
rect 179266 706522 179502 706758
rect 179586 706522 179822 706758
rect 179266 706202 179502 706438
rect 179586 706202 179822 706438
rect 179266 690658 179502 690894
rect 179586 690658 179822 690894
rect 179266 690338 179502 690574
rect 179586 690338 179822 690574
rect 179266 656658 179502 656894
rect 179586 656658 179822 656894
rect 179266 656338 179502 656574
rect 179586 656338 179822 656574
rect 179266 622658 179502 622894
rect 179586 622658 179822 622894
rect 179266 622338 179502 622574
rect 179586 622338 179822 622574
rect 179266 588658 179502 588894
rect 179586 588658 179822 588894
rect 179266 588338 179502 588574
rect 179586 588338 179822 588574
rect 179266 554658 179502 554894
rect 179586 554658 179822 554894
rect 179266 554338 179502 554574
rect 179586 554338 179822 554574
rect 179266 520658 179502 520894
rect 179586 520658 179822 520894
rect 179266 520338 179502 520574
rect 179586 520338 179822 520574
rect 179266 486658 179502 486894
rect 179586 486658 179822 486894
rect 179266 486338 179502 486574
rect 179586 486338 179822 486574
rect 179266 452658 179502 452894
rect 179586 452658 179822 452894
rect 179266 452338 179502 452574
rect 179586 452338 179822 452574
rect 179266 418658 179502 418894
rect 179586 418658 179822 418894
rect 179266 418338 179502 418574
rect 179586 418338 179822 418574
rect 179266 384658 179502 384894
rect 179586 384658 179822 384894
rect 179266 384338 179502 384574
rect 179586 384338 179822 384574
rect 179266 350658 179502 350894
rect 179586 350658 179822 350894
rect 179266 350338 179502 350574
rect 179586 350338 179822 350574
rect 179266 316658 179502 316894
rect 179586 316658 179822 316894
rect 179266 316338 179502 316574
rect 179586 316338 179822 316574
rect 179266 282658 179502 282894
rect 179586 282658 179822 282894
rect 179266 282338 179502 282574
rect 179586 282338 179822 282574
rect 179266 248658 179502 248894
rect 179586 248658 179822 248894
rect 179266 248338 179502 248574
rect 179586 248338 179822 248574
rect 182986 707482 183222 707718
rect 183306 707482 183542 707718
rect 182986 707162 183222 707398
rect 183306 707162 183542 707398
rect 182986 694378 183222 694614
rect 183306 694378 183542 694614
rect 182986 694058 183222 694294
rect 183306 694058 183542 694294
rect 182986 660378 183222 660614
rect 183306 660378 183542 660614
rect 182986 660058 183222 660294
rect 183306 660058 183542 660294
rect 182986 626378 183222 626614
rect 183306 626378 183542 626614
rect 182986 626058 183222 626294
rect 183306 626058 183542 626294
rect 182986 592378 183222 592614
rect 183306 592378 183542 592614
rect 182986 592058 183222 592294
rect 183306 592058 183542 592294
rect 182986 558378 183222 558614
rect 183306 558378 183542 558614
rect 182986 558058 183222 558294
rect 183306 558058 183542 558294
rect 182986 524378 183222 524614
rect 183306 524378 183542 524614
rect 182986 524058 183222 524294
rect 183306 524058 183542 524294
rect 182986 490378 183222 490614
rect 183306 490378 183542 490614
rect 182986 490058 183222 490294
rect 183306 490058 183542 490294
rect 182986 456378 183222 456614
rect 183306 456378 183542 456614
rect 182986 456058 183222 456294
rect 183306 456058 183542 456294
rect 182986 422378 183222 422614
rect 183306 422378 183542 422614
rect 182986 422058 183222 422294
rect 183306 422058 183542 422294
rect 182986 388378 183222 388614
rect 183306 388378 183542 388614
rect 182986 388058 183222 388294
rect 183306 388058 183542 388294
rect 182986 354378 183222 354614
rect 183306 354378 183542 354614
rect 182986 354058 183222 354294
rect 183306 354058 183542 354294
rect 182986 320378 183222 320614
rect 183306 320378 183542 320614
rect 182986 320058 183222 320294
rect 183306 320058 183542 320294
rect 182986 286378 183222 286614
rect 183306 286378 183542 286614
rect 182986 286058 183222 286294
rect 183306 286058 183542 286294
rect 182986 252378 183222 252614
rect 183306 252378 183542 252614
rect 182986 252058 183222 252294
rect 183306 252058 183542 252294
rect 186706 708442 186942 708678
rect 187026 708442 187262 708678
rect 186706 708122 186942 708358
rect 187026 708122 187262 708358
rect 186706 698098 186942 698334
rect 187026 698098 187262 698334
rect 186706 697778 186942 698014
rect 187026 697778 187262 698014
rect 186706 664098 186942 664334
rect 187026 664098 187262 664334
rect 186706 663778 186942 664014
rect 187026 663778 187262 664014
rect 186706 630098 186942 630334
rect 187026 630098 187262 630334
rect 186706 629778 186942 630014
rect 187026 629778 187262 630014
rect 186706 596098 186942 596334
rect 187026 596098 187262 596334
rect 186706 595778 186942 596014
rect 187026 595778 187262 596014
rect 186706 562098 186942 562334
rect 187026 562098 187262 562334
rect 186706 561778 186942 562014
rect 187026 561778 187262 562014
rect 186706 528098 186942 528334
rect 187026 528098 187262 528334
rect 186706 527778 186942 528014
rect 187026 527778 187262 528014
rect 186706 494098 186942 494334
rect 187026 494098 187262 494334
rect 186706 493778 186942 494014
rect 187026 493778 187262 494014
rect 186706 460098 186942 460334
rect 187026 460098 187262 460334
rect 186706 459778 186942 460014
rect 187026 459778 187262 460014
rect 186706 426098 186942 426334
rect 187026 426098 187262 426334
rect 186706 425778 186942 426014
rect 187026 425778 187262 426014
rect 186706 392098 186942 392334
rect 187026 392098 187262 392334
rect 186706 391778 186942 392014
rect 187026 391778 187262 392014
rect 186706 358098 186942 358334
rect 187026 358098 187262 358334
rect 186706 357778 186942 358014
rect 187026 357778 187262 358014
rect 186706 324098 186942 324334
rect 187026 324098 187262 324334
rect 186706 323778 186942 324014
rect 187026 323778 187262 324014
rect 186706 290098 186942 290334
rect 187026 290098 187262 290334
rect 186706 289778 186942 290014
rect 187026 289778 187262 290014
rect 186706 256098 186942 256334
rect 187026 256098 187262 256334
rect 186706 255778 186942 256014
rect 187026 255778 187262 256014
rect 190426 709402 190662 709638
rect 190746 709402 190982 709638
rect 190426 709082 190662 709318
rect 190746 709082 190982 709318
rect 190426 667818 190662 668054
rect 190746 667818 190982 668054
rect 190426 667498 190662 667734
rect 190746 667498 190982 667734
rect 190426 633818 190662 634054
rect 190746 633818 190982 634054
rect 190426 633498 190662 633734
rect 190746 633498 190982 633734
rect 190426 599818 190662 600054
rect 190746 599818 190982 600054
rect 190426 599498 190662 599734
rect 190746 599498 190982 599734
rect 190426 565818 190662 566054
rect 190746 565818 190982 566054
rect 190426 565498 190662 565734
rect 190746 565498 190982 565734
rect 190426 531818 190662 532054
rect 190746 531818 190982 532054
rect 190426 531498 190662 531734
rect 190746 531498 190982 531734
rect 190426 497818 190662 498054
rect 190746 497818 190982 498054
rect 190426 497498 190662 497734
rect 190746 497498 190982 497734
rect 190426 463818 190662 464054
rect 190746 463818 190982 464054
rect 190426 463498 190662 463734
rect 190746 463498 190982 463734
rect 190426 429818 190662 430054
rect 190746 429818 190982 430054
rect 190426 429498 190662 429734
rect 190746 429498 190982 429734
rect 190426 395818 190662 396054
rect 190746 395818 190982 396054
rect 190426 395498 190662 395734
rect 190746 395498 190982 395734
rect 190426 361818 190662 362054
rect 190746 361818 190982 362054
rect 190426 361498 190662 361734
rect 190746 361498 190982 361734
rect 190426 327818 190662 328054
rect 190746 327818 190982 328054
rect 190426 327498 190662 327734
rect 190746 327498 190982 327734
rect 190426 293818 190662 294054
rect 190746 293818 190982 294054
rect 190426 293498 190662 293734
rect 190746 293498 190982 293734
rect 190426 259818 190662 260054
rect 190746 259818 190982 260054
rect 190426 259498 190662 259734
rect 190746 259498 190982 259734
rect 190426 225818 190662 226054
rect 190746 225818 190982 226054
rect 190426 225498 190662 225734
rect 190746 225498 190982 225734
rect 194146 710362 194382 710598
rect 194466 710362 194702 710598
rect 194146 710042 194382 710278
rect 194466 710042 194702 710278
rect 194146 671538 194382 671774
rect 194466 671538 194702 671774
rect 194146 671218 194382 671454
rect 194466 671218 194702 671454
rect 194146 637538 194382 637774
rect 194466 637538 194702 637774
rect 194146 637218 194382 637454
rect 194466 637218 194702 637454
rect 194146 603538 194382 603774
rect 194466 603538 194702 603774
rect 194146 603218 194382 603454
rect 194466 603218 194702 603454
rect 194146 569538 194382 569774
rect 194466 569538 194702 569774
rect 194146 569218 194382 569454
rect 194466 569218 194702 569454
rect 194146 535538 194382 535774
rect 194466 535538 194702 535774
rect 194146 535218 194382 535454
rect 194466 535218 194702 535454
rect 194146 501538 194382 501774
rect 194466 501538 194702 501774
rect 194146 501218 194382 501454
rect 194466 501218 194702 501454
rect 194146 467538 194382 467774
rect 194466 467538 194702 467774
rect 194146 467218 194382 467454
rect 194466 467218 194702 467454
rect 194146 433538 194382 433774
rect 194466 433538 194702 433774
rect 194146 433218 194382 433454
rect 194466 433218 194702 433454
rect 194146 399538 194382 399774
rect 194466 399538 194702 399774
rect 194146 399218 194382 399454
rect 194466 399218 194702 399454
rect 194146 365538 194382 365774
rect 194466 365538 194702 365774
rect 194146 365218 194382 365454
rect 194466 365218 194702 365454
rect 194146 331538 194382 331774
rect 194466 331538 194702 331774
rect 194146 331218 194382 331454
rect 194466 331218 194702 331454
rect 194146 297538 194382 297774
rect 194466 297538 194702 297774
rect 194146 297218 194382 297454
rect 194466 297218 194702 297454
rect 194146 263538 194382 263774
rect 194466 263538 194702 263774
rect 194146 263218 194382 263454
rect 194466 263218 194702 263454
rect 194146 229538 194382 229774
rect 194466 229538 194702 229774
rect 194146 229218 194382 229454
rect 194466 229218 194702 229454
rect 197866 711322 198102 711558
rect 198186 711322 198422 711558
rect 197866 711002 198102 711238
rect 198186 711002 198422 711238
rect 197866 675258 198102 675494
rect 198186 675258 198422 675494
rect 197866 674938 198102 675174
rect 198186 674938 198422 675174
rect 197866 641258 198102 641494
rect 198186 641258 198422 641494
rect 197866 640938 198102 641174
rect 198186 640938 198422 641174
rect 197866 607258 198102 607494
rect 198186 607258 198422 607494
rect 197866 606938 198102 607174
rect 198186 606938 198422 607174
rect 197866 573258 198102 573494
rect 198186 573258 198422 573494
rect 197866 572938 198102 573174
rect 198186 572938 198422 573174
rect 197866 539258 198102 539494
rect 198186 539258 198422 539494
rect 197866 538938 198102 539174
rect 198186 538938 198422 539174
rect 197866 505258 198102 505494
rect 198186 505258 198422 505494
rect 197866 504938 198102 505174
rect 198186 504938 198422 505174
rect 197866 471258 198102 471494
rect 198186 471258 198422 471494
rect 197866 470938 198102 471174
rect 198186 470938 198422 471174
rect 197866 437258 198102 437494
rect 198186 437258 198422 437494
rect 197866 436938 198102 437174
rect 198186 436938 198422 437174
rect 197866 403258 198102 403494
rect 198186 403258 198422 403494
rect 197866 402938 198102 403174
rect 198186 402938 198422 403174
rect 197866 369258 198102 369494
rect 198186 369258 198422 369494
rect 197866 368938 198102 369174
rect 198186 368938 198422 369174
rect 197866 335258 198102 335494
rect 198186 335258 198422 335494
rect 197866 334938 198102 335174
rect 198186 334938 198422 335174
rect 197866 301258 198102 301494
rect 198186 301258 198422 301494
rect 197866 300938 198102 301174
rect 198186 300938 198422 301174
rect 197866 267258 198102 267494
rect 198186 267258 198422 267494
rect 197866 266938 198102 267174
rect 198186 266938 198422 267174
rect 197866 233258 198102 233494
rect 198186 233258 198422 233494
rect 197866 232938 198102 233174
rect 198186 232938 198422 233174
rect 205826 704602 206062 704838
rect 206146 704602 206382 704838
rect 205826 704282 206062 704518
rect 206146 704282 206382 704518
rect 205826 683218 206062 683454
rect 206146 683218 206382 683454
rect 205826 682898 206062 683134
rect 206146 682898 206382 683134
rect 205826 649218 206062 649454
rect 206146 649218 206382 649454
rect 205826 648898 206062 649134
rect 206146 648898 206382 649134
rect 205826 615218 206062 615454
rect 206146 615218 206382 615454
rect 205826 614898 206062 615134
rect 206146 614898 206382 615134
rect 205826 581218 206062 581454
rect 206146 581218 206382 581454
rect 205826 580898 206062 581134
rect 206146 580898 206382 581134
rect 205826 547218 206062 547454
rect 206146 547218 206382 547454
rect 205826 546898 206062 547134
rect 206146 546898 206382 547134
rect 205826 513218 206062 513454
rect 206146 513218 206382 513454
rect 205826 512898 206062 513134
rect 206146 512898 206382 513134
rect 205826 479218 206062 479454
rect 206146 479218 206382 479454
rect 205826 478898 206062 479134
rect 206146 478898 206382 479134
rect 205826 445218 206062 445454
rect 206146 445218 206382 445454
rect 205826 444898 206062 445134
rect 206146 444898 206382 445134
rect 205826 411218 206062 411454
rect 206146 411218 206382 411454
rect 205826 410898 206062 411134
rect 206146 410898 206382 411134
rect 205826 377218 206062 377454
rect 206146 377218 206382 377454
rect 205826 376898 206062 377134
rect 206146 376898 206382 377134
rect 205826 343218 206062 343454
rect 206146 343218 206382 343454
rect 205826 342898 206062 343134
rect 206146 342898 206382 343134
rect 205826 309218 206062 309454
rect 206146 309218 206382 309454
rect 205826 308898 206062 309134
rect 206146 308898 206382 309134
rect 205826 275218 206062 275454
rect 206146 275218 206382 275454
rect 205826 274898 206062 275134
rect 206146 274898 206382 275134
rect 205826 241218 206062 241454
rect 206146 241218 206382 241454
rect 205826 240898 206062 241134
rect 206146 240898 206382 241134
rect 209546 705562 209782 705798
rect 209866 705562 210102 705798
rect 209546 705242 209782 705478
rect 209866 705242 210102 705478
rect 209546 686938 209782 687174
rect 209866 686938 210102 687174
rect 209546 686618 209782 686854
rect 209866 686618 210102 686854
rect 209546 652938 209782 653174
rect 209866 652938 210102 653174
rect 209546 652618 209782 652854
rect 209866 652618 210102 652854
rect 209546 618938 209782 619174
rect 209866 618938 210102 619174
rect 209546 618618 209782 618854
rect 209866 618618 210102 618854
rect 209546 584938 209782 585174
rect 209866 584938 210102 585174
rect 209546 584618 209782 584854
rect 209866 584618 210102 584854
rect 209546 550938 209782 551174
rect 209866 550938 210102 551174
rect 209546 550618 209782 550854
rect 209866 550618 210102 550854
rect 209546 516938 209782 517174
rect 209866 516938 210102 517174
rect 209546 516618 209782 516854
rect 209866 516618 210102 516854
rect 209546 482938 209782 483174
rect 209866 482938 210102 483174
rect 209546 482618 209782 482854
rect 209866 482618 210102 482854
rect 209546 448938 209782 449174
rect 209866 448938 210102 449174
rect 209546 448618 209782 448854
rect 209866 448618 210102 448854
rect 209546 414938 209782 415174
rect 209866 414938 210102 415174
rect 209546 414618 209782 414854
rect 209866 414618 210102 414854
rect 209546 380938 209782 381174
rect 209866 380938 210102 381174
rect 209546 380618 209782 380854
rect 209866 380618 210102 380854
rect 209546 346938 209782 347174
rect 209866 346938 210102 347174
rect 209546 346618 209782 346854
rect 209866 346618 210102 346854
rect 209546 312938 209782 313174
rect 209866 312938 210102 313174
rect 209546 312618 209782 312854
rect 209866 312618 210102 312854
rect 209546 278938 209782 279174
rect 209866 278938 210102 279174
rect 209546 278618 209782 278854
rect 209866 278618 210102 278854
rect 209546 244938 209782 245174
rect 209866 244938 210102 245174
rect 209546 244618 209782 244854
rect 209866 244618 210102 244854
rect 213266 706522 213502 706758
rect 213586 706522 213822 706758
rect 213266 706202 213502 706438
rect 213586 706202 213822 706438
rect 213266 690658 213502 690894
rect 213586 690658 213822 690894
rect 213266 690338 213502 690574
rect 213586 690338 213822 690574
rect 213266 656658 213502 656894
rect 213586 656658 213822 656894
rect 213266 656338 213502 656574
rect 213586 656338 213822 656574
rect 213266 622658 213502 622894
rect 213586 622658 213822 622894
rect 213266 622338 213502 622574
rect 213586 622338 213822 622574
rect 213266 588658 213502 588894
rect 213586 588658 213822 588894
rect 213266 588338 213502 588574
rect 213586 588338 213822 588574
rect 213266 554658 213502 554894
rect 213586 554658 213822 554894
rect 213266 554338 213502 554574
rect 213586 554338 213822 554574
rect 213266 520658 213502 520894
rect 213586 520658 213822 520894
rect 213266 520338 213502 520574
rect 213586 520338 213822 520574
rect 213266 486658 213502 486894
rect 213586 486658 213822 486894
rect 213266 486338 213502 486574
rect 213586 486338 213822 486574
rect 213266 452658 213502 452894
rect 213586 452658 213822 452894
rect 213266 452338 213502 452574
rect 213586 452338 213822 452574
rect 213266 418658 213502 418894
rect 213586 418658 213822 418894
rect 213266 418338 213502 418574
rect 213586 418338 213822 418574
rect 213266 384658 213502 384894
rect 213586 384658 213822 384894
rect 213266 384338 213502 384574
rect 213586 384338 213822 384574
rect 213266 350658 213502 350894
rect 213586 350658 213822 350894
rect 213266 350338 213502 350574
rect 213586 350338 213822 350574
rect 213266 316658 213502 316894
rect 213586 316658 213822 316894
rect 213266 316338 213502 316574
rect 213586 316338 213822 316574
rect 213266 282658 213502 282894
rect 213586 282658 213822 282894
rect 213266 282338 213502 282574
rect 213586 282338 213822 282574
rect 213266 248658 213502 248894
rect 213586 248658 213822 248894
rect 213266 248338 213502 248574
rect 213586 248338 213822 248574
rect 216986 707482 217222 707718
rect 217306 707482 217542 707718
rect 216986 707162 217222 707398
rect 217306 707162 217542 707398
rect 216986 694378 217222 694614
rect 217306 694378 217542 694614
rect 216986 694058 217222 694294
rect 217306 694058 217542 694294
rect 216986 660378 217222 660614
rect 217306 660378 217542 660614
rect 216986 660058 217222 660294
rect 217306 660058 217542 660294
rect 216986 626378 217222 626614
rect 217306 626378 217542 626614
rect 216986 626058 217222 626294
rect 217306 626058 217542 626294
rect 216986 592378 217222 592614
rect 217306 592378 217542 592614
rect 216986 592058 217222 592294
rect 217306 592058 217542 592294
rect 216986 558378 217222 558614
rect 217306 558378 217542 558614
rect 216986 558058 217222 558294
rect 217306 558058 217542 558294
rect 216986 524378 217222 524614
rect 217306 524378 217542 524614
rect 216986 524058 217222 524294
rect 217306 524058 217542 524294
rect 216986 490378 217222 490614
rect 217306 490378 217542 490614
rect 216986 490058 217222 490294
rect 217306 490058 217542 490294
rect 216986 456378 217222 456614
rect 217306 456378 217542 456614
rect 216986 456058 217222 456294
rect 217306 456058 217542 456294
rect 216986 422378 217222 422614
rect 217306 422378 217542 422614
rect 216986 422058 217222 422294
rect 217306 422058 217542 422294
rect 216986 388378 217222 388614
rect 217306 388378 217542 388614
rect 216986 388058 217222 388294
rect 217306 388058 217542 388294
rect 216986 354378 217222 354614
rect 217306 354378 217542 354614
rect 216986 354058 217222 354294
rect 217306 354058 217542 354294
rect 216986 320378 217222 320614
rect 217306 320378 217542 320614
rect 216986 320058 217222 320294
rect 217306 320058 217542 320294
rect 216986 286378 217222 286614
rect 217306 286378 217542 286614
rect 216986 286058 217222 286294
rect 217306 286058 217542 286294
rect 216986 252378 217222 252614
rect 217306 252378 217542 252614
rect 216986 252058 217222 252294
rect 217306 252058 217542 252294
rect 220706 708442 220942 708678
rect 221026 708442 221262 708678
rect 220706 708122 220942 708358
rect 221026 708122 221262 708358
rect 220706 698098 220942 698334
rect 221026 698098 221262 698334
rect 220706 697778 220942 698014
rect 221026 697778 221262 698014
rect 220706 664098 220942 664334
rect 221026 664098 221262 664334
rect 220706 663778 220942 664014
rect 221026 663778 221262 664014
rect 220706 630098 220942 630334
rect 221026 630098 221262 630334
rect 220706 629778 220942 630014
rect 221026 629778 221262 630014
rect 220706 596098 220942 596334
rect 221026 596098 221262 596334
rect 220706 595778 220942 596014
rect 221026 595778 221262 596014
rect 220706 562098 220942 562334
rect 221026 562098 221262 562334
rect 220706 561778 220942 562014
rect 221026 561778 221262 562014
rect 220706 528098 220942 528334
rect 221026 528098 221262 528334
rect 220706 527778 220942 528014
rect 221026 527778 221262 528014
rect 220706 494098 220942 494334
rect 221026 494098 221262 494334
rect 220706 493778 220942 494014
rect 221026 493778 221262 494014
rect 220706 460098 220942 460334
rect 221026 460098 221262 460334
rect 220706 459778 220942 460014
rect 221026 459778 221262 460014
rect 220706 426098 220942 426334
rect 221026 426098 221262 426334
rect 220706 425778 220942 426014
rect 221026 425778 221262 426014
rect 220706 392098 220942 392334
rect 221026 392098 221262 392334
rect 220706 391778 220942 392014
rect 221026 391778 221262 392014
rect 220706 358098 220942 358334
rect 221026 358098 221262 358334
rect 220706 357778 220942 358014
rect 221026 357778 221262 358014
rect 220706 324098 220942 324334
rect 221026 324098 221262 324334
rect 220706 323778 220942 324014
rect 221026 323778 221262 324014
rect 220706 290098 220942 290334
rect 221026 290098 221262 290334
rect 220706 289778 220942 290014
rect 221026 289778 221262 290014
rect 220706 256098 220942 256334
rect 221026 256098 221262 256334
rect 220706 255778 220942 256014
rect 221026 255778 221262 256014
rect 160146 195538 160382 195774
rect 160466 195538 160702 195774
rect 160146 195218 160382 195454
rect 160466 195218 160702 195454
rect 163866 199258 164102 199494
rect 164186 199258 164422 199494
rect 163866 198938 164102 199174
rect 164186 198938 164422 199174
rect 134376 188098 134612 188334
rect 134696 188098 134932 188334
rect 135016 188098 135252 188334
rect 135336 188098 135572 188334
rect 135656 188098 135892 188334
rect 135976 188098 136212 188334
rect 136296 188098 136532 188334
rect 136616 188098 136852 188334
rect 136936 188098 137172 188334
rect 137256 188098 137492 188334
rect 137576 188098 137812 188334
rect 137896 188098 138132 188334
rect 138216 188098 138452 188334
rect 138536 188098 138772 188334
rect 138856 188098 139092 188334
rect 139176 188098 139412 188334
rect 139496 188098 139732 188334
rect 139816 188098 140052 188334
rect 140136 188098 140372 188334
rect 140456 188098 140692 188334
rect 140776 188098 141012 188334
rect 141096 188098 141332 188334
rect 141416 188098 141652 188334
rect 141736 188098 141972 188334
rect 142056 188098 142292 188334
rect 142376 188098 142612 188334
rect 142696 188098 142932 188334
rect 143016 188098 143252 188334
rect 143336 188098 143572 188334
rect 143656 188098 143892 188334
rect 143976 188098 144212 188334
rect 144296 188098 144532 188334
rect 144616 188098 144852 188334
rect 144936 188098 145172 188334
rect 145256 188098 145492 188334
rect 145576 188098 145812 188334
rect 145896 188098 146132 188334
rect 146216 188098 146452 188334
rect 146536 188098 146772 188334
rect 146856 188098 147092 188334
rect 147176 188098 147412 188334
rect 147496 188098 147732 188334
rect 147816 188098 148052 188334
rect 148136 188098 148372 188334
rect 148456 188098 148692 188334
rect 148776 188098 149012 188334
rect 149096 188098 149332 188334
rect 149416 188098 149652 188334
rect 149736 188098 149972 188334
rect 150056 188098 150292 188334
rect 150376 188098 150612 188334
rect 150696 188098 150932 188334
rect 151016 188098 151252 188334
rect 151336 188098 151572 188334
rect 151656 188098 151892 188334
rect 151976 188098 152212 188334
rect 152296 188098 152532 188334
rect 152616 188098 152852 188334
rect 152936 188098 153172 188334
rect 153256 188098 153492 188334
rect 153576 188098 153812 188334
rect 153896 188098 154132 188334
rect 154216 188098 154452 188334
rect 154536 188098 154772 188334
rect 154856 188098 155092 188334
rect 155176 188098 155412 188334
rect 155496 188098 155732 188334
rect 155816 188098 156052 188334
rect 156136 188098 156372 188334
rect 156456 188098 156692 188334
rect 156776 188098 157012 188334
rect 157096 188098 157332 188334
rect 157416 188098 157652 188334
rect 157736 188098 157972 188334
rect 158056 188098 158292 188334
rect 158376 188098 158612 188334
rect 158696 188098 158932 188334
rect 159016 188098 159252 188334
rect 159336 188098 159572 188334
rect 159656 188098 159892 188334
rect 159976 188098 160212 188334
rect 160296 188098 160532 188334
rect 160616 188098 160852 188334
rect 160936 188098 161172 188334
rect 161256 188098 161492 188334
rect 161576 188098 161812 188334
rect 161896 188098 162132 188334
rect 162216 188098 162452 188334
rect 134376 187778 134612 188014
rect 134696 187778 134932 188014
rect 135016 187778 135252 188014
rect 135336 187778 135572 188014
rect 135656 187778 135892 188014
rect 135976 187778 136212 188014
rect 136296 187778 136532 188014
rect 136616 187778 136852 188014
rect 136936 187778 137172 188014
rect 137256 187778 137492 188014
rect 137576 187778 137812 188014
rect 137896 187778 138132 188014
rect 138216 187778 138452 188014
rect 138536 187778 138772 188014
rect 138856 187778 139092 188014
rect 139176 187778 139412 188014
rect 139496 187778 139732 188014
rect 139816 187778 140052 188014
rect 140136 187778 140372 188014
rect 140456 187778 140692 188014
rect 140776 187778 141012 188014
rect 141096 187778 141332 188014
rect 141416 187778 141652 188014
rect 141736 187778 141972 188014
rect 142056 187778 142292 188014
rect 142376 187778 142612 188014
rect 142696 187778 142932 188014
rect 143016 187778 143252 188014
rect 143336 187778 143572 188014
rect 143656 187778 143892 188014
rect 143976 187778 144212 188014
rect 144296 187778 144532 188014
rect 144616 187778 144852 188014
rect 144936 187778 145172 188014
rect 145256 187778 145492 188014
rect 145576 187778 145812 188014
rect 145896 187778 146132 188014
rect 146216 187778 146452 188014
rect 146536 187778 146772 188014
rect 146856 187778 147092 188014
rect 147176 187778 147412 188014
rect 147496 187778 147732 188014
rect 147816 187778 148052 188014
rect 148136 187778 148372 188014
rect 148456 187778 148692 188014
rect 148776 187778 149012 188014
rect 149096 187778 149332 188014
rect 149416 187778 149652 188014
rect 149736 187778 149972 188014
rect 150056 187778 150292 188014
rect 150376 187778 150612 188014
rect 150696 187778 150932 188014
rect 151016 187778 151252 188014
rect 151336 187778 151572 188014
rect 151656 187778 151892 188014
rect 151976 187778 152212 188014
rect 152296 187778 152532 188014
rect 152616 187778 152852 188014
rect 152936 187778 153172 188014
rect 153256 187778 153492 188014
rect 153576 187778 153812 188014
rect 153896 187778 154132 188014
rect 154216 187778 154452 188014
rect 154536 187778 154772 188014
rect 154856 187778 155092 188014
rect 155176 187778 155412 188014
rect 155496 187778 155732 188014
rect 155816 187778 156052 188014
rect 156136 187778 156372 188014
rect 156456 187778 156692 188014
rect 156776 187778 157012 188014
rect 157096 187778 157332 188014
rect 157416 187778 157652 188014
rect 157736 187778 157972 188014
rect 158056 187778 158292 188014
rect 158376 187778 158612 188014
rect 158696 187778 158932 188014
rect 159016 187778 159252 188014
rect 159336 187778 159572 188014
rect 159656 187778 159892 188014
rect 159976 187778 160212 188014
rect 160296 187778 160532 188014
rect 160616 187778 160852 188014
rect 160936 187778 161172 188014
rect 161256 187778 161492 188014
rect 161576 187778 161812 188014
rect 161896 187778 162132 188014
rect 162216 187778 162452 188014
rect 129866 165258 130102 165494
rect 130186 165258 130422 165494
rect 129866 164938 130102 165174
rect 130186 164938 130422 165174
rect 134446 161545 134682 161781
rect 134766 161545 135002 161781
rect 145266 180658 145502 180894
rect 145586 180658 145822 180894
rect 145266 180338 145502 180574
rect 145586 180338 145822 180574
rect 148986 184378 149222 184614
rect 149306 184378 149542 184614
rect 148986 184058 149222 184294
rect 149306 184058 149542 184294
rect 137826 173218 138062 173454
rect 138146 173218 138382 173454
rect 137826 172898 138062 173134
rect 138146 172898 138382 173134
rect 134446 161225 134682 161461
rect 134766 161225 135002 161461
rect 160146 161538 160382 161774
rect 160466 161538 160702 161774
rect 160146 161218 160382 161454
rect 160466 161218 160702 161454
rect 163866 165258 164102 165494
rect 164186 165258 164422 165494
rect 163866 164938 164102 165174
rect 164186 164938 164422 165174
rect 171826 207218 172062 207454
rect 172146 207218 172382 207454
rect 171826 206898 172062 207134
rect 172146 206898 172382 207134
rect 171826 173218 172062 173454
rect 172146 173218 172382 173454
rect 171826 172898 172062 173134
rect 172146 172898 172382 173134
rect 171826 139218 172062 139454
rect 172146 139218 172382 139454
rect 171826 138898 172062 139134
rect 172146 138898 172382 139134
rect 114986 116378 115222 116614
rect 115306 116378 115542 116614
rect 114986 116058 115222 116294
rect 115306 116058 115542 116294
rect 135610 108938 135846 109174
rect 135610 108618 135846 108854
rect 166330 108938 166566 109174
rect 166330 108618 166566 108854
rect 120250 105218 120486 105454
rect 120250 104898 120486 105134
rect 150970 105218 151206 105454
rect 150970 104898 151206 105134
rect 171826 105218 172062 105454
rect 172146 105218 172382 105454
rect 171826 104898 172062 105134
rect 172146 104898 172382 105134
rect 114986 82378 115222 82614
rect 115306 82378 115542 82614
rect 114986 82058 115222 82294
rect 115306 82058 115542 82294
rect 114986 48378 115222 48614
rect 115306 48378 115542 48614
rect 114986 48058 115222 48294
rect 115306 48058 115542 48294
rect 114986 14378 115222 14614
rect 115306 14378 115542 14614
rect 114986 14058 115222 14294
rect 115306 14058 115542 14294
rect 114986 -3462 115222 -3226
rect 115306 -3462 115542 -3226
rect 114986 -3782 115222 -3546
rect 115306 -3782 115542 -3546
rect 118706 52098 118942 52334
rect 119026 52098 119262 52334
rect 118706 51778 118942 52014
rect 119026 51778 119262 52014
rect 118706 18098 118942 18334
rect 119026 18098 119262 18334
rect 118706 17778 118942 18014
rect 119026 17778 119262 18014
rect 118706 -4422 118942 -4186
rect 119026 -4422 119262 -4186
rect 118706 -4742 118942 -4506
rect 119026 -4742 119262 -4506
rect 122426 55818 122662 56054
rect 122746 55818 122982 56054
rect 122426 55498 122662 55734
rect 122746 55498 122982 55734
rect 126146 59538 126382 59774
rect 126466 59538 126702 59774
rect 126146 59218 126382 59454
rect 126466 59218 126702 59454
rect 122426 21818 122662 22054
rect 122746 21818 122982 22054
rect 122426 21498 122662 21734
rect 122746 21498 122982 21734
rect 122426 -5382 122662 -5146
rect 122746 -5382 122982 -5146
rect 122426 -5702 122662 -5466
rect 122746 -5702 122982 -5466
rect 126146 25538 126382 25774
rect 126466 25538 126702 25774
rect 126146 25218 126382 25454
rect 126466 25218 126702 25454
rect 129866 63258 130102 63494
rect 130186 63258 130422 63494
rect 129866 62938 130102 63174
rect 130186 62938 130422 63174
rect 129866 29258 130102 29494
rect 130186 29258 130422 29494
rect 129866 28938 130102 29174
rect 130186 28938 130422 29174
rect 126146 -6342 126382 -6106
rect 126466 -6342 126702 -6106
rect 126146 -6662 126382 -6426
rect 126466 -6662 126702 -6426
rect 137826 71218 138062 71454
rect 138146 71218 138382 71454
rect 137826 70898 138062 71134
rect 138146 70898 138382 71134
rect 137826 37218 138062 37454
rect 138146 37218 138382 37454
rect 137826 36898 138062 37134
rect 138146 36898 138382 37134
rect 141546 40938 141782 41174
rect 141866 40938 142102 41174
rect 141546 40618 141782 40854
rect 141866 40618 142102 40854
rect 141546 6938 141782 7174
rect 141866 6938 142102 7174
rect 141546 6618 141782 6854
rect 141866 6618 142102 6854
rect 129866 -7302 130102 -7066
rect 130186 -7302 130422 -7066
rect 129866 -7622 130102 -7386
rect 130186 -7622 130422 -7386
rect 137826 3218 138062 3454
rect 138146 3218 138382 3454
rect 137826 2898 138062 3134
rect 138146 2898 138382 3134
rect 137826 -582 138062 -346
rect 138146 -582 138382 -346
rect 137826 -902 138062 -666
rect 138146 -902 138382 -666
rect 145266 44658 145502 44894
rect 145586 44658 145822 44894
rect 145266 44338 145502 44574
rect 145586 44338 145822 44574
rect 145266 10658 145502 10894
rect 145586 10658 145822 10894
rect 145266 10338 145502 10574
rect 145586 10338 145822 10574
rect 141546 -1542 141782 -1306
rect 141866 -1542 142102 -1306
rect 141546 -1862 141782 -1626
rect 141866 -1862 142102 -1626
rect 148986 48378 149222 48614
rect 149306 48378 149542 48614
rect 148986 48058 149222 48294
rect 149306 48058 149542 48294
rect 148986 14378 149222 14614
rect 149306 14378 149542 14614
rect 148986 14058 149222 14294
rect 149306 14058 149542 14294
rect 145266 -2502 145502 -2266
rect 145586 -2502 145822 -2266
rect 145266 -2822 145502 -2586
rect 145586 -2822 145822 -2586
rect 152706 52098 152942 52334
rect 153026 52098 153262 52334
rect 152706 51778 152942 52014
rect 153026 51778 153262 52014
rect 152706 18098 152942 18334
rect 153026 18098 153262 18334
rect 152706 17778 152942 18014
rect 153026 17778 153262 18014
rect 148986 -3462 149222 -3226
rect 149306 -3462 149542 -3226
rect 148986 -3782 149222 -3546
rect 149306 -3782 149542 -3546
rect 156426 55818 156662 56054
rect 156746 55818 156982 56054
rect 156426 55498 156662 55734
rect 156746 55498 156982 55734
rect 156426 21818 156662 22054
rect 156746 21818 156982 22054
rect 156426 21498 156662 21734
rect 156746 21498 156982 21734
rect 152706 -4422 152942 -4186
rect 153026 -4422 153262 -4186
rect 152706 -4742 152942 -4506
rect 153026 -4742 153262 -4506
rect 160146 59538 160382 59774
rect 160466 59538 160702 59774
rect 160146 59218 160382 59454
rect 160466 59218 160702 59454
rect 160146 25538 160382 25774
rect 160466 25538 160702 25774
rect 160146 25218 160382 25454
rect 160466 25218 160702 25454
rect 156426 -5382 156662 -5146
rect 156746 -5382 156982 -5146
rect 156426 -5702 156662 -5466
rect 156746 -5702 156982 -5466
rect 163866 63258 164102 63494
rect 164186 63258 164422 63494
rect 163866 62938 164102 63174
rect 164186 62938 164422 63174
rect 163866 29258 164102 29494
rect 164186 29258 164422 29494
rect 163866 28938 164102 29174
rect 164186 28938 164422 29174
rect 160146 -6342 160382 -6106
rect 160466 -6342 160702 -6106
rect 160146 -6662 160382 -6426
rect 160466 -6662 160702 -6426
rect 171826 71218 172062 71454
rect 172146 71218 172382 71454
rect 171826 70898 172062 71134
rect 172146 70898 172382 71134
rect 171826 37218 172062 37454
rect 172146 37218 172382 37454
rect 171826 36898 172062 37134
rect 172146 36898 172382 37134
rect 163866 -7302 164102 -7066
rect 164186 -7302 164422 -7066
rect 163866 -7622 164102 -7386
rect 164186 -7622 164422 -7386
rect 171826 3218 172062 3454
rect 172146 3218 172382 3454
rect 171826 2898 172062 3134
rect 172146 2898 172382 3134
rect 171826 -582 172062 -346
rect 172146 -582 172382 -346
rect 171826 -902 172062 -666
rect 172146 -902 172382 -666
rect 175546 210938 175782 211174
rect 175866 210938 176102 211174
rect 175546 210618 175782 210854
rect 175866 210618 176102 210854
rect 175546 176938 175782 177174
rect 175866 176938 176102 177174
rect 175546 176618 175782 176854
rect 175866 176618 176102 176854
rect 175546 142938 175782 143174
rect 175866 142938 176102 143174
rect 175546 142618 175782 142854
rect 175866 142618 176102 142854
rect 175546 108938 175782 109174
rect 175866 108938 176102 109174
rect 175546 108618 175782 108854
rect 175866 108618 176102 108854
rect 175546 74938 175782 75174
rect 175866 74938 176102 75174
rect 175546 74618 175782 74854
rect 175866 74618 176102 74854
rect 175546 40938 175782 41174
rect 175866 40938 176102 41174
rect 175546 40618 175782 40854
rect 175866 40618 176102 40854
rect 175546 6938 175782 7174
rect 175866 6938 176102 7174
rect 175546 6618 175782 6854
rect 175866 6618 176102 6854
rect 175546 -1542 175782 -1306
rect 175866 -1542 176102 -1306
rect 175546 -1862 175782 -1626
rect 175866 -1862 176102 -1626
rect 179266 180658 179502 180894
rect 179586 180658 179822 180894
rect 179266 180338 179502 180574
rect 179586 180338 179822 180574
rect 179266 146658 179502 146894
rect 179586 146658 179822 146894
rect 179266 146338 179502 146574
rect 179586 146338 179822 146574
rect 179266 112658 179502 112894
rect 179586 112658 179822 112894
rect 179266 112338 179502 112574
rect 179586 112338 179822 112574
rect 179266 78658 179502 78894
rect 179586 78658 179822 78894
rect 179266 78338 179502 78574
rect 179586 78338 179822 78574
rect 179266 44658 179502 44894
rect 179586 44658 179822 44894
rect 179266 44338 179502 44574
rect 179586 44338 179822 44574
rect 179266 10658 179502 10894
rect 179586 10658 179822 10894
rect 179266 10338 179502 10574
rect 179586 10338 179822 10574
rect 179266 -2502 179502 -2266
rect 179586 -2502 179822 -2266
rect 179266 -2822 179502 -2586
rect 179586 -2822 179822 -2586
rect 182986 184378 183222 184614
rect 183306 184378 183542 184614
rect 182986 184058 183222 184294
rect 183306 184058 183542 184294
rect 182986 150378 183222 150614
rect 183306 150378 183542 150614
rect 182986 150058 183222 150294
rect 183306 150058 183542 150294
rect 182986 116378 183222 116614
rect 183306 116378 183542 116614
rect 182986 116058 183222 116294
rect 183306 116058 183542 116294
rect 182986 82378 183222 82614
rect 183306 82378 183542 82614
rect 182986 82058 183222 82294
rect 183306 82058 183542 82294
rect 182986 48378 183222 48614
rect 183306 48378 183542 48614
rect 182986 48058 183222 48294
rect 183306 48058 183542 48294
rect 182986 14378 183222 14614
rect 183306 14378 183542 14614
rect 182986 14058 183222 14294
rect 183306 14058 183542 14294
rect 182986 -3462 183222 -3226
rect 183306 -3462 183542 -3226
rect 182986 -3782 183222 -3546
rect 183306 -3782 183542 -3546
rect 186706 188098 186942 188334
rect 187026 188098 187262 188334
rect 186706 187778 186942 188014
rect 187026 187778 187262 188014
rect 186706 154098 186942 154334
rect 187026 154098 187262 154334
rect 186706 153778 186942 154014
rect 187026 153778 187262 154014
rect 186706 120098 186942 120334
rect 187026 120098 187262 120334
rect 186706 119778 186942 120014
rect 187026 119778 187262 120014
rect 186706 86098 186942 86334
rect 187026 86098 187262 86334
rect 186706 85778 186942 86014
rect 187026 85778 187262 86014
rect 186706 52098 186942 52334
rect 187026 52098 187262 52334
rect 186706 51778 186942 52014
rect 187026 51778 187262 52014
rect 186706 18098 186942 18334
rect 187026 18098 187262 18334
rect 186706 17778 186942 18014
rect 187026 17778 187262 18014
rect 186706 -4422 186942 -4186
rect 187026 -4422 187262 -4186
rect 186706 -4742 186942 -4506
rect 187026 -4742 187262 -4506
rect 224426 709402 224662 709638
rect 224746 709402 224982 709638
rect 224426 709082 224662 709318
rect 224746 709082 224982 709318
rect 224426 667818 224662 668054
rect 224746 667818 224982 668054
rect 224426 667498 224662 667734
rect 224746 667498 224982 667734
rect 224426 633818 224662 634054
rect 224746 633818 224982 634054
rect 224426 633498 224662 633734
rect 224746 633498 224982 633734
rect 224426 599818 224662 600054
rect 224746 599818 224982 600054
rect 224426 599498 224662 599734
rect 224746 599498 224982 599734
rect 224426 565818 224662 566054
rect 224746 565818 224982 566054
rect 224426 565498 224662 565734
rect 224746 565498 224982 565734
rect 224426 531818 224662 532054
rect 224746 531818 224982 532054
rect 224426 531498 224662 531734
rect 224746 531498 224982 531734
rect 224426 497818 224662 498054
rect 224746 497818 224982 498054
rect 224426 497498 224662 497734
rect 224746 497498 224982 497734
rect 224426 463818 224662 464054
rect 224746 463818 224982 464054
rect 224426 463498 224662 463734
rect 224746 463498 224982 463734
rect 224426 429818 224662 430054
rect 224746 429818 224982 430054
rect 224426 429498 224662 429734
rect 224746 429498 224982 429734
rect 224426 395818 224662 396054
rect 224746 395818 224982 396054
rect 224426 395498 224662 395734
rect 224746 395498 224982 395734
rect 224426 361818 224662 362054
rect 224746 361818 224982 362054
rect 224426 361498 224662 361734
rect 224746 361498 224982 361734
rect 224426 327818 224662 328054
rect 224746 327818 224982 328054
rect 224426 327498 224662 327734
rect 224746 327498 224982 327734
rect 224426 293818 224662 294054
rect 224746 293818 224982 294054
rect 224426 293498 224662 293734
rect 224746 293498 224982 293734
rect 224426 259818 224662 260054
rect 224746 259818 224982 260054
rect 224426 259498 224662 259734
rect 224746 259498 224982 259734
rect 224426 225755 224662 225991
rect 224746 225755 224982 225991
rect 228146 710362 228382 710598
rect 228466 710362 228702 710598
rect 228146 710042 228382 710278
rect 228466 710042 228702 710278
rect 228146 671538 228382 671774
rect 228466 671538 228702 671774
rect 228146 671218 228382 671454
rect 228466 671218 228702 671454
rect 228146 637538 228382 637774
rect 228466 637538 228702 637774
rect 228146 637218 228382 637454
rect 228466 637218 228702 637454
rect 228146 603538 228382 603774
rect 228466 603538 228702 603774
rect 228146 603218 228382 603454
rect 228466 603218 228702 603454
rect 228146 569538 228382 569774
rect 228466 569538 228702 569774
rect 228146 569218 228382 569454
rect 228466 569218 228702 569454
rect 228146 535538 228382 535774
rect 228466 535538 228702 535774
rect 228146 535218 228382 535454
rect 228466 535218 228702 535454
rect 228146 501538 228382 501774
rect 228466 501538 228702 501774
rect 228146 501218 228382 501454
rect 228466 501218 228702 501454
rect 228146 467538 228382 467774
rect 228466 467538 228702 467774
rect 228146 467218 228382 467454
rect 228466 467218 228702 467454
rect 228146 433538 228382 433774
rect 228466 433538 228702 433774
rect 228146 433218 228382 433454
rect 228466 433218 228702 433454
rect 228146 399538 228382 399774
rect 228466 399538 228702 399774
rect 228146 399218 228382 399454
rect 228466 399218 228702 399454
rect 228146 365538 228382 365774
rect 228466 365538 228702 365774
rect 228146 365218 228382 365454
rect 228466 365218 228702 365454
rect 228146 331538 228382 331774
rect 228466 331538 228702 331774
rect 228146 331218 228382 331454
rect 228466 331218 228702 331454
rect 228146 297538 228382 297774
rect 228466 297538 228702 297774
rect 228146 297218 228382 297454
rect 228466 297218 228702 297454
rect 228146 263538 228382 263774
rect 228466 263538 228702 263774
rect 228146 263218 228382 263454
rect 228466 263218 228702 263454
rect 228146 229538 228382 229774
rect 228466 229538 228702 229774
rect 228146 229218 228382 229454
rect 228466 229218 228702 229454
rect 231866 711322 232102 711558
rect 232186 711322 232422 711558
rect 231866 711002 232102 711238
rect 232186 711002 232422 711238
rect 231866 675258 232102 675494
rect 232186 675258 232422 675494
rect 231866 674938 232102 675174
rect 232186 674938 232422 675174
rect 231866 641258 232102 641494
rect 232186 641258 232422 641494
rect 231866 640938 232102 641174
rect 232186 640938 232422 641174
rect 231866 607258 232102 607494
rect 232186 607258 232422 607494
rect 231866 606938 232102 607174
rect 232186 606938 232422 607174
rect 231866 573258 232102 573494
rect 232186 573258 232422 573494
rect 231866 572938 232102 573174
rect 232186 572938 232422 573174
rect 231866 539258 232102 539494
rect 232186 539258 232422 539494
rect 231866 538938 232102 539174
rect 232186 538938 232422 539174
rect 231866 505258 232102 505494
rect 232186 505258 232422 505494
rect 231866 504938 232102 505174
rect 232186 504938 232422 505174
rect 231866 471258 232102 471494
rect 232186 471258 232422 471494
rect 231866 470938 232102 471174
rect 232186 470938 232422 471174
rect 231866 437258 232102 437494
rect 232186 437258 232422 437494
rect 231866 436938 232102 437174
rect 232186 436938 232422 437174
rect 231866 403258 232102 403494
rect 232186 403258 232422 403494
rect 231866 402938 232102 403174
rect 232186 402938 232422 403174
rect 231866 369258 232102 369494
rect 232186 369258 232422 369494
rect 231866 368938 232102 369174
rect 232186 368938 232422 369174
rect 231866 335258 232102 335494
rect 232186 335258 232422 335494
rect 231866 334938 232102 335174
rect 232186 334938 232422 335174
rect 231866 301258 232102 301494
rect 232186 301258 232422 301494
rect 231866 300938 232102 301174
rect 232186 300938 232422 301174
rect 231866 267258 232102 267494
rect 232186 267258 232422 267494
rect 231866 266938 232102 267174
rect 232186 266938 232422 267174
rect 231866 233258 232102 233494
rect 232186 233258 232422 233494
rect 231866 232938 232102 233174
rect 232186 232938 232422 233174
rect 239826 704602 240062 704838
rect 240146 704602 240382 704838
rect 239826 704282 240062 704518
rect 240146 704282 240382 704518
rect 239826 683218 240062 683454
rect 240146 683218 240382 683454
rect 239826 682898 240062 683134
rect 240146 682898 240382 683134
rect 239826 649218 240062 649454
rect 240146 649218 240382 649454
rect 239826 648898 240062 649134
rect 240146 648898 240382 649134
rect 239826 615218 240062 615454
rect 240146 615218 240382 615454
rect 239826 614898 240062 615134
rect 240146 614898 240382 615134
rect 239826 581218 240062 581454
rect 240146 581218 240382 581454
rect 239826 580898 240062 581134
rect 240146 580898 240382 581134
rect 239826 547218 240062 547454
rect 240146 547218 240382 547454
rect 239826 546898 240062 547134
rect 240146 546898 240382 547134
rect 239826 513218 240062 513454
rect 240146 513218 240382 513454
rect 239826 512898 240062 513134
rect 240146 512898 240382 513134
rect 239826 479218 240062 479454
rect 240146 479218 240382 479454
rect 239826 478898 240062 479134
rect 240146 478898 240382 479134
rect 239826 445218 240062 445454
rect 240146 445218 240382 445454
rect 239826 444898 240062 445134
rect 240146 444898 240382 445134
rect 239826 411218 240062 411454
rect 240146 411218 240382 411454
rect 239826 410898 240062 411134
rect 240146 410898 240382 411134
rect 239826 377218 240062 377454
rect 240146 377218 240382 377454
rect 239826 376898 240062 377134
rect 240146 376898 240382 377134
rect 239826 343218 240062 343454
rect 240146 343218 240382 343454
rect 239826 342898 240062 343134
rect 240146 342898 240382 343134
rect 239826 309218 240062 309454
rect 240146 309218 240382 309454
rect 239826 308898 240062 309134
rect 240146 308898 240382 309134
rect 239826 275218 240062 275454
rect 240146 275218 240382 275454
rect 239826 274898 240062 275134
rect 240146 274898 240382 275134
rect 239826 241218 240062 241454
rect 240146 241218 240382 241454
rect 239826 240898 240062 241134
rect 240146 240898 240382 241134
rect 243546 705562 243782 705798
rect 243866 705562 244102 705798
rect 243546 705242 243782 705478
rect 243866 705242 244102 705478
rect 243546 686938 243782 687174
rect 243866 686938 244102 687174
rect 243546 686618 243782 686854
rect 243866 686618 244102 686854
rect 243546 652938 243782 653174
rect 243866 652938 244102 653174
rect 243546 652618 243782 652854
rect 243866 652618 244102 652854
rect 243546 618938 243782 619174
rect 243866 618938 244102 619174
rect 243546 618618 243782 618854
rect 243866 618618 244102 618854
rect 243546 584938 243782 585174
rect 243866 584938 244102 585174
rect 243546 584618 243782 584854
rect 243866 584618 244102 584854
rect 243546 550938 243782 551174
rect 243866 550938 244102 551174
rect 243546 550618 243782 550854
rect 243866 550618 244102 550854
rect 243546 516938 243782 517174
rect 243866 516938 244102 517174
rect 243546 516618 243782 516854
rect 243866 516618 244102 516854
rect 243546 482938 243782 483174
rect 243866 482938 244102 483174
rect 243546 482618 243782 482854
rect 243866 482618 244102 482854
rect 243546 448938 243782 449174
rect 243866 448938 244102 449174
rect 243546 448618 243782 448854
rect 243866 448618 244102 448854
rect 243546 414938 243782 415174
rect 243866 414938 244102 415174
rect 243546 414618 243782 414854
rect 243866 414618 244102 414854
rect 243546 380938 243782 381174
rect 243866 380938 244102 381174
rect 243546 380618 243782 380854
rect 243866 380618 244102 380854
rect 243546 346938 243782 347174
rect 243866 346938 244102 347174
rect 243546 346618 243782 346854
rect 243866 346618 244102 346854
rect 243546 312938 243782 313174
rect 243866 312938 244102 313174
rect 243546 312618 243782 312854
rect 243866 312618 244102 312854
rect 243546 278938 243782 279174
rect 243866 278938 244102 279174
rect 243546 278618 243782 278854
rect 243866 278618 244102 278854
rect 243546 244938 243782 245174
rect 243866 244938 244102 245174
rect 243546 244618 243782 244854
rect 243866 244618 244102 244854
rect 247266 706522 247502 706758
rect 247586 706522 247822 706758
rect 247266 706202 247502 706438
rect 247586 706202 247822 706438
rect 247266 690658 247502 690894
rect 247586 690658 247822 690894
rect 247266 690338 247502 690574
rect 247586 690338 247822 690574
rect 247266 656658 247502 656894
rect 247586 656658 247822 656894
rect 247266 656338 247502 656574
rect 247586 656338 247822 656574
rect 247266 622658 247502 622894
rect 247586 622658 247822 622894
rect 247266 622338 247502 622574
rect 247586 622338 247822 622574
rect 247266 588658 247502 588894
rect 247586 588658 247822 588894
rect 247266 588338 247502 588574
rect 247586 588338 247822 588574
rect 247266 554658 247502 554894
rect 247586 554658 247822 554894
rect 247266 554338 247502 554574
rect 247586 554338 247822 554574
rect 247266 520658 247502 520894
rect 247586 520658 247822 520894
rect 247266 520338 247502 520574
rect 247586 520338 247822 520574
rect 247266 486658 247502 486894
rect 247586 486658 247822 486894
rect 247266 486338 247502 486574
rect 247586 486338 247822 486574
rect 247266 452658 247502 452894
rect 247586 452658 247822 452894
rect 247266 452338 247502 452574
rect 247586 452338 247822 452574
rect 247266 418658 247502 418894
rect 247586 418658 247822 418894
rect 247266 418338 247502 418574
rect 247586 418338 247822 418574
rect 247266 384658 247502 384894
rect 247586 384658 247822 384894
rect 247266 384338 247502 384574
rect 247586 384338 247822 384574
rect 247266 350658 247502 350894
rect 247586 350658 247822 350894
rect 247266 350338 247502 350574
rect 247586 350338 247822 350574
rect 247266 316658 247502 316894
rect 247586 316658 247822 316894
rect 247266 316338 247502 316574
rect 247586 316338 247822 316574
rect 247266 282658 247502 282894
rect 247586 282658 247822 282894
rect 247266 282338 247502 282574
rect 247586 282338 247822 282574
rect 247266 248658 247502 248894
rect 247586 248658 247822 248894
rect 247266 248338 247502 248574
rect 247586 248338 247822 248574
rect 250986 707482 251222 707718
rect 251306 707482 251542 707718
rect 250986 707162 251222 707398
rect 251306 707162 251542 707398
rect 250986 694378 251222 694614
rect 251306 694378 251542 694614
rect 250986 694058 251222 694294
rect 251306 694058 251542 694294
rect 250986 660378 251222 660614
rect 251306 660378 251542 660614
rect 250986 660058 251222 660294
rect 251306 660058 251542 660294
rect 250986 626378 251222 626614
rect 251306 626378 251542 626614
rect 250986 626058 251222 626294
rect 251306 626058 251542 626294
rect 250986 592378 251222 592614
rect 251306 592378 251542 592614
rect 250986 592058 251222 592294
rect 251306 592058 251542 592294
rect 250986 558378 251222 558614
rect 251306 558378 251542 558614
rect 250986 558058 251222 558294
rect 251306 558058 251542 558294
rect 250986 524378 251222 524614
rect 251306 524378 251542 524614
rect 250986 524058 251222 524294
rect 251306 524058 251542 524294
rect 250986 490378 251222 490614
rect 251306 490378 251542 490614
rect 250986 490058 251222 490294
rect 251306 490058 251542 490294
rect 250986 456378 251222 456614
rect 251306 456378 251542 456614
rect 250986 456058 251222 456294
rect 251306 456058 251542 456294
rect 250986 422378 251222 422614
rect 251306 422378 251542 422614
rect 250986 422058 251222 422294
rect 251306 422058 251542 422294
rect 250986 388378 251222 388614
rect 251306 388378 251542 388614
rect 250986 388058 251222 388294
rect 251306 388058 251542 388294
rect 250986 354378 251222 354614
rect 251306 354378 251542 354614
rect 250986 354058 251222 354294
rect 251306 354058 251542 354294
rect 250986 320378 251222 320614
rect 251306 320378 251542 320614
rect 250986 320058 251222 320294
rect 251306 320058 251542 320294
rect 250986 286378 251222 286614
rect 251306 286378 251542 286614
rect 250986 286058 251222 286294
rect 251306 286058 251542 286294
rect 250986 252378 251222 252614
rect 251306 252378 251542 252614
rect 250986 252058 251222 252294
rect 251306 252058 251542 252294
rect 220706 222098 220942 222334
rect 221026 222098 221262 222334
rect 220706 221778 220942 222014
rect 221026 221778 221262 222014
rect 190426 191818 190662 192054
rect 190746 191818 190982 192054
rect 190426 191498 190662 191734
rect 190746 191498 190982 191734
rect 190426 157818 190662 158054
rect 190746 157818 190982 158054
rect 190426 157498 190662 157734
rect 190746 157498 190982 157734
rect 190426 123818 190662 124054
rect 190746 123818 190982 124054
rect 190426 123498 190662 123734
rect 190746 123498 190982 123734
rect 190426 89818 190662 90054
rect 190746 89818 190982 90054
rect 190426 89498 190662 89734
rect 190746 89498 190982 89734
rect 190426 55818 190662 56054
rect 190746 55818 190982 56054
rect 190426 55498 190662 55734
rect 190746 55498 190982 55734
rect 190426 21818 190662 22054
rect 190746 21818 190982 22054
rect 190426 21498 190662 21734
rect 190746 21498 190982 21734
rect 190426 -5382 190662 -5146
rect 190746 -5382 190982 -5146
rect 190426 -5702 190662 -5466
rect 190746 -5702 190982 -5466
rect 194146 195538 194382 195774
rect 194466 195538 194702 195774
rect 194146 195218 194382 195454
rect 194466 195218 194702 195454
rect 194146 161538 194382 161774
rect 194466 161538 194702 161774
rect 194146 161218 194382 161454
rect 194466 161218 194702 161454
rect 194146 127538 194382 127774
rect 194466 127538 194702 127774
rect 194146 127218 194382 127454
rect 194466 127218 194702 127454
rect 194146 93538 194382 93774
rect 194466 93538 194702 93774
rect 194146 93218 194382 93454
rect 194466 93218 194702 93454
rect 194146 59538 194382 59774
rect 194466 59538 194702 59774
rect 194146 59218 194382 59454
rect 194466 59218 194702 59454
rect 194146 25538 194382 25774
rect 194466 25538 194702 25774
rect 194146 25218 194382 25454
rect 194466 25218 194702 25454
rect 194146 -6342 194382 -6106
rect 194466 -6342 194702 -6106
rect 194146 -6662 194382 -6426
rect 194466 -6662 194702 -6426
rect 197866 199258 198102 199494
rect 198186 199258 198422 199494
rect 197866 198938 198102 199174
rect 198186 198938 198422 199174
rect 197866 165258 198102 165494
rect 198186 165258 198422 165494
rect 197866 164938 198102 165174
rect 198186 164938 198422 165174
rect 197866 131258 198102 131494
rect 198186 131258 198422 131494
rect 197866 130938 198102 131174
rect 198186 130938 198422 131174
rect 197866 97258 198102 97494
rect 198186 97258 198422 97494
rect 197866 96938 198102 97174
rect 198186 96938 198422 97174
rect 197866 63258 198102 63494
rect 198186 63258 198422 63494
rect 197866 62938 198102 63174
rect 198186 62938 198422 63174
rect 197866 29258 198102 29494
rect 198186 29258 198422 29494
rect 197866 28938 198102 29174
rect 198186 28938 198422 29174
rect 197866 -7302 198102 -7066
rect 198186 -7302 198422 -7066
rect 197866 -7622 198102 -7386
rect 198186 -7622 198422 -7386
rect 205826 207218 206062 207454
rect 206146 207218 206382 207454
rect 205826 206898 206062 207134
rect 206146 206898 206382 207134
rect 205826 173218 206062 173454
rect 206146 173218 206382 173454
rect 205826 172898 206062 173134
rect 206146 172898 206382 173134
rect 205826 139218 206062 139454
rect 206146 139218 206382 139454
rect 205826 138898 206062 139134
rect 206146 138898 206382 139134
rect 205826 105218 206062 105454
rect 206146 105218 206382 105454
rect 205826 104898 206062 105134
rect 206146 104898 206382 105134
rect 205826 71218 206062 71454
rect 206146 71218 206382 71454
rect 205826 70898 206062 71134
rect 206146 70898 206382 71134
rect 205826 37218 206062 37454
rect 206146 37218 206382 37454
rect 205826 36898 206062 37134
rect 206146 36898 206382 37134
rect 205826 3218 206062 3454
rect 206146 3218 206382 3454
rect 205826 2898 206062 3134
rect 206146 2898 206382 3134
rect 205826 -582 206062 -346
rect 206146 -582 206382 -346
rect 205826 -902 206062 -666
rect 206146 -902 206382 -666
rect 209546 210938 209782 211174
rect 209866 210938 210102 211174
rect 209546 210618 209782 210854
rect 209866 210618 210102 210854
rect 209546 176938 209782 177174
rect 209866 176938 210102 177174
rect 209546 176618 209782 176854
rect 209866 176618 210102 176854
rect 209546 142938 209782 143174
rect 209866 142938 210102 143174
rect 209546 142618 209782 142854
rect 209866 142618 210102 142854
rect 209546 108938 209782 109174
rect 209866 108938 210102 109174
rect 209546 108618 209782 108854
rect 209866 108618 210102 108854
rect 209546 74938 209782 75174
rect 209866 74938 210102 75174
rect 209546 74618 209782 74854
rect 209866 74618 210102 74854
rect 209546 40938 209782 41174
rect 209866 40938 210102 41174
rect 209546 40618 209782 40854
rect 209866 40618 210102 40854
rect 209546 6938 209782 7174
rect 209866 6938 210102 7174
rect 209546 6618 209782 6854
rect 209866 6618 210102 6854
rect 209546 -1542 209782 -1306
rect 209866 -1542 210102 -1306
rect 209546 -1862 209782 -1626
rect 209866 -1862 210102 -1626
rect 213266 180658 213502 180894
rect 213586 180658 213822 180894
rect 213266 180338 213502 180574
rect 213586 180338 213822 180574
rect 213266 146658 213502 146894
rect 213586 146658 213822 146894
rect 213266 146338 213502 146574
rect 213586 146338 213822 146574
rect 213266 112658 213502 112894
rect 213586 112658 213822 112894
rect 213266 112338 213502 112574
rect 213586 112338 213822 112574
rect 213266 78658 213502 78894
rect 213586 78658 213822 78894
rect 213266 78338 213502 78574
rect 213586 78338 213822 78574
rect 213266 44658 213502 44894
rect 213586 44658 213822 44894
rect 213266 44338 213502 44574
rect 213586 44338 213822 44574
rect 213266 10658 213502 10894
rect 213586 10658 213822 10894
rect 213266 10338 213502 10574
rect 213586 10338 213822 10574
rect 213266 -2502 213502 -2266
rect 213586 -2502 213822 -2266
rect 213266 -2822 213502 -2586
rect 213586 -2822 213822 -2586
rect 216986 184378 217222 184614
rect 217306 184378 217542 184614
rect 216986 184058 217222 184294
rect 217306 184058 217542 184294
rect 216986 150378 217222 150614
rect 217306 150378 217542 150614
rect 216986 150058 217222 150294
rect 217306 150058 217542 150294
rect 216986 116378 217222 116614
rect 217306 116378 217542 116614
rect 216986 116058 217222 116294
rect 217306 116058 217542 116294
rect 216986 82378 217222 82614
rect 217306 82378 217542 82614
rect 216986 82058 217222 82294
rect 217306 82058 217542 82294
rect 216986 48378 217222 48614
rect 217306 48378 217542 48614
rect 216986 48058 217222 48294
rect 217306 48058 217542 48294
rect 216986 14378 217222 14614
rect 217306 14378 217542 14614
rect 216986 14058 217222 14294
rect 217306 14058 217542 14294
rect 216986 -3462 217222 -3226
rect 217306 -3462 217542 -3226
rect 216986 -3782 217222 -3546
rect 217306 -3782 217542 -3546
rect 254706 708442 254942 708678
rect 255026 708442 255262 708678
rect 254706 708122 254942 708358
rect 255026 708122 255262 708358
rect 254706 698098 254942 698334
rect 255026 698098 255262 698334
rect 254706 697778 254942 698014
rect 255026 697778 255262 698014
rect 254706 664098 254942 664334
rect 255026 664098 255262 664334
rect 254706 663778 254942 664014
rect 255026 663778 255262 664014
rect 254706 630098 254942 630334
rect 255026 630098 255262 630334
rect 254706 629778 254942 630014
rect 255026 629778 255262 630014
rect 254706 596098 254942 596334
rect 255026 596098 255262 596334
rect 254706 595778 254942 596014
rect 255026 595778 255262 596014
rect 254706 562098 254942 562334
rect 255026 562098 255262 562334
rect 254706 561778 254942 562014
rect 255026 561778 255262 562014
rect 254706 528098 254942 528334
rect 255026 528098 255262 528334
rect 254706 527778 254942 528014
rect 255026 527778 255262 528014
rect 254706 494098 254942 494334
rect 255026 494098 255262 494334
rect 254706 493778 254942 494014
rect 255026 493778 255262 494014
rect 254706 460098 254942 460334
rect 255026 460098 255262 460334
rect 254706 459778 254942 460014
rect 255026 459778 255262 460014
rect 254706 426098 254942 426334
rect 255026 426098 255262 426334
rect 254706 425778 254942 426014
rect 255026 425778 255262 426014
rect 254706 392098 254942 392334
rect 255026 392098 255262 392334
rect 254706 391778 254942 392014
rect 255026 391778 255262 392014
rect 254706 358098 254942 358334
rect 255026 358098 255262 358334
rect 254706 357778 254942 358014
rect 255026 357778 255262 358014
rect 254706 324098 254942 324334
rect 255026 324098 255262 324334
rect 254706 323778 254942 324014
rect 255026 323778 255262 324014
rect 254706 290098 254942 290334
rect 255026 290098 255262 290334
rect 254706 289778 254942 290014
rect 255026 289778 255262 290014
rect 254706 256098 254942 256334
rect 255026 256098 255262 256334
rect 254706 255778 254942 256014
rect 255026 255778 255262 256014
rect 258426 709402 258662 709638
rect 258746 709402 258982 709638
rect 258426 709082 258662 709318
rect 258746 709082 258982 709318
rect 258426 667818 258662 668054
rect 258746 667818 258982 668054
rect 258426 667498 258662 667734
rect 258746 667498 258982 667734
rect 258426 633818 258662 634054
rect 258746 633818 258982 634054
rect 258426 633498 258662 633734
rect 258746 633498 258982 633734
rect 258426 599818 258662 600054
rect 258746 599818 258982 600054
rect 258426 599498 258662 599734
rect 258746 599498 258982 599734
rect 258426 565818 258662 566054
rect 258746 565818 258982 566054
rect 258426 565498 258662 565734
rect 258746 565498 258982 565734
rect 258426 531818 258662 532054
rect 258746 531818 258982 532054
rect 258426 531498 258662 531734
rect 258746 531498 258982 531734
rect 258426 497818 258662 498054
rect 258746 497818 258982 498054
rect 258426 497498 258662 497734
rect 258746 497498 258982 497734
rect 258426 463818 258662 464054
rect 258746 463818 258982 464054
rect 258426 463498 258662 463734
rect 258746 463498 258982 463734
rect 258426 429818 258662 430054
rect 258746 429818 258982 430054
rect 258426 429498 258662 429734
rect 258746 429498 258982 429734
rect 258426 395818 258662 396054
rect 258746 395818 258982 396054
rect 258426 395498 258662 395734
rect 258746 395498 258982 395734
rect 258426 361818 258662 362054
rect 258746 361818 258982 362054
rect 258426 361498 258662 361734
rect 258746 361498 258982 361734
rect 258426 327818 258662 328054
rect 258746 327818 258982 328054
rect 258426 327498 258662 327734
rect 258746 327498 258982 327734
rect 258426 293818 258662 294054
rect 258746 293818 258982 294054
rect 258426 293498 258662 293734
rect 258746 293498 258982 293734
rect 258426 259818 258662 260054
rect 258746 259818 258982 260054
rect 258426 259498 258662 259734
rect 258746 259498 258982 259734
rect 258426 225755 258662 225991
rect 258746 225755 258982 225991
rect 262146 710362 262382 710598
rect 262466 710362 262702 710598
rect 262146 710042 262382 710278
rect 262466 710042 262702 710278
rect 262146 671538 262382 671774
rect 262466 671538 262702 671774
rect 262146 671218 262382 671454
rect 262466 671218 262702 671454
rect 262146 637538 262382 637774
rect 262466 637538 262702 637774
rect 262146 637218 262382 637454
rect 262466 637218 262702 637454
rect 262146 603538 262382 603774
rect 262466 603538 262702 603774
rect 262146 603218 262382 603454
rect 262466 603218 262702 603454
rect 262146 569538 262382 569774
rect 262466 569538 262702 569774
rect 262146 569218 262382 569454
rect 262466 569218 262702 569454
rect 262146 535538 262382 535774
rect 262466 535538 262702 535774
rect 262146 535218 262382 535454
rect 262466 535218 262702 535454
rect 262146 501538 262382 501774
rect 262466 501538 262702 501774
rect 262146 501218 262382 501454
rect 262466 501218 262702 501454
rect 262146 467538 262382 467774
rect 262466 467538 262702 467774
rect 262146 467218 262382 467454
rect 262466 467218 262702 467454
rect 262146 433538 262382 433774
rect 262466 433538 262702 433774
rect 262146 433218 262382 433454
rect 262466 433218 262702 433454
rect 262146 399538 262382 399774
rect 262466 399538 262702 399774
rect 262146 399218 262382 399454
rect 262466 399218 262702 399454
rect 262146 365538 262382 365774
rect 262466 365538 262702 365774
rect 262146 365218 262382 365454
rect 262466 365218 262702 365454
rect 262146 331538 262382 331774
rect 262466 331538 262702 331774
rect 262146 331218 262382 331454
rect 262466 331218 262702 331454
rect 262146 297538 262382 297774
rect 262466 297538 262702 297774
rect 262146 297218 262382 297454
rect 262466 297218 262702 297454
rect 262146 263538 262382 263774
rect 262466 263538 262702 263774
rect 262146 263218 262382 263454
rect 262466 263218 262702 263454
rect 262146 229538 262382 229774
rect 262466 229538 262702 229774
rect 262146 229218 262382 229454
rect 262466 229218 262702 229454
rect 265866 711322 266102 711558
rect 266186 711322 266422 711558
rect 265866 711002 266102 711238
rect 266186 711002 266422 711238
rect 265866 675258 266102 675494
rect 266186 675258 266422 675494
rect 265866 674938 266102 675174
rect 266186 674938 266422 675174
rect 265866 641258 266102 641494
rect 266186 641258 266422 641494
rect 265866 640938 266102 641174
rect 266186 640938 266422 641174
rect 265866 607258 266102 607494
rect 266186 607258 266422 607494
rect 265866 606938 266102 607174
rect 266186 606938 266422 607174
rect 265866 573258 266102 573494
rect 266186 573258 266422 573494
rect 265866 572938 266102 573174
rect 266186 572938 266422 573174
rect 265866 539258 266102 539494
rect 266186 539258 266422 539494
rect 265866 538938 266102 539174
rect 266186 538938 266422 539174
rect 265866 505258 266102 505494
rect 266186 505258 266422 505494
rect 265866 504938 266102 505174
rect 266186 504938 266422 505174
rect 265866 471258 266102 471494
rect 266186 471258 266422 471494
rect 265866 470938 266102 471174
rect 266186 470938 266422 471174
rect 265866 437258 266102 437494
rect 266186 437258 266422 437494
rect 265866 436938 266102 437174
rect 266186 436938 266422 437174
rect 265866 403258 266102 403494
rect 266186 403258 266422 403494
rect 265866 402938 266102 403174
rect 266186 402938 266422 403174
rect 265866 369258 266102 369494
rect 266186 369258 266422 369494
rect 265866 368938 266102 369174
rect 266186 368938 266422 369174
rect 265866 335258 266102 335494
rect 266186 335258 266422 335494
rect 265866 334938 266102 335174
rect 266186 334938 266422 335174
rect 265866 301258 266102 301494
rect 266186 301258 266422 301494
rect 265866 300938 266102 301174
rect 266186 300938 266422 301174
rect 265866 267258 266102 267494
rect 266186 267258 266422 267494
rect 265866 266938 266102 267174
rect 266186 266938 266422 267174
rect 265866 233258 266102 233494
rect 266186 233258 266422 233494
rect 265866 232938 266102 233174
rect 266186 232938 266422 233174
rect 273826 704602 274062 704838
rect 274146 704602 274382 704838
rect 273826 704282 274062 704518
rect 274146 704282 274382 704518
rect 273826 683218 274062 683454
rect 274146 683218 274382 683454
rect 273826 682898 274062 683134
rect 274146 682898 274382 683134
rect 273826 649218 274062 649454
rect 274146 649218 274382 649454
rect 273826 648898 274062 649134
rect 274146 648898 274382 649134
rect 273826 615218 274062 615454
rect 274146 615218 274382 615454
rect 273826 614898 274062 615134
rect 274146 614898 274382 615134
rect 273826 581218 274062 581454
rect 274146 581218 274382 581454
rect 273826 580898 274062 581134
rect 274146 580898 274382 581134
rect 273826 547218 274062 547454
rect 274146 547218 274382 547454
rect 273826 546898 274062 547134
rect 274146 546898 274382 547134
rect 273826 513218 274062 513454
rect 274146 513218 274382 513454
rect 273826 512898 274062 513134
rect 274146 512898 274382 513134
rect 273826 479218 274062 479454
rect 274146 479218 274382 479454
rect 273826 478898 274062 479134
rect 274146 478898 274382 479134
rect 273826 445218 274062 445454
rect 274146 445218 274382 445454
rect 273826 444898 274062 445134
rect 274146 444898 274382 445134
rect 273826 411218 274062 411454
rect 274146 411218 274382 411454
rect 273826 410898 274062 411134
rect 274146 410898 274382 411134
rect 273826 377218 274062 377454
rect 274146 377218 274382 377454
rect 273826 376898 274062 377134
rect 274146 376898 274382 377134
rect 273826 343218 274062 343454
rect 274146 343218 274382 343454
rect 273826 342898 274062 343134
rect 274146 342898 274382 343134
rect 273826 309218 274062 309454
rect 274146 309218 274382 309454
rect 273826 308898 274062 309134
rect 274146 308898 274382 309134
rect 273826 275218 274062 275454
rect 274146 275218 274382 275454
rect 273826 274898 274062 275134
rect 274146 274898 274382 275134
rect 273826 241218 274062 241454
rect 274146 241218 274382 241454
rect 273826 240898 274062 241134
rect 274146 240898 274382 241134
rect 277546 705562 277782 705798
rect 277866 705562 278102 705798
rect 277546 705242 277782 705478
rect 277866 705242 278102 705478
rect 277546 686938 277782 687174
rect 277866 686938 278102 687174
rect 277546 686618 277782 686854
rect 277866 686618 278102 686854
rect 277546 652938 277782 653174
rect 277866 652938 278102 653174
rect 277546 652618 277782 652854
rect 277866 652618 278102 652854
rect 277546 618938 277782 619174
rect 277866 618938 278102 619174
rect 277546 618618 277782 618854
rect 277866 618618 278102 618854
rect 277546 584938 277782 585174
rect 277866 584938 278102 585174
rect 277546 584618 277782 584854
rect 277866 584618 278102 584854
rect 277546 550938 277782 551174
rect 277866 550938 278102 551174
rect 277546 550618 277782 550854
rect 277866 550618 278102 550854
rect 277546 516938 277782 517174
rect 277866 516938 278102 517174
rect 277546 516618 277782 516854
rect 277866 516618 278102 516854
rect 277546 482938 277782 483174
rect 277866 482938 278102 483174
rect 277546 482618 277782 482854
rect 277866 482618 278102 482854
rect 277546 448938 277782 449174
rect 277866 448938 278102 449174
rect 277546 448618 277782 448854
rect 277866 448618 278102 448854
rect 277546 414938 277782 415174
rect 277866 414938 278102 415174
rect 277546 414618 277782 414854
rect 277866 414618 278102 414854
rect 277546 380938 277782 381174
rect 277866 380938 278102 381174
rect 277546 380618 277782 380854
rect 277866 380618 278102 380854
rect 277546 346938 277782 347174
rect 277866 346938 278102 347174
rect 277546 346618 277782 346854
rect 277866 346618 278102 346854
rect 277546 312938 277782 313174
rect 277866 312938 278102 313174
rect 277546 312618 277782 312854
rect 277866 312618 278102 312854
rect 277546 278938 277782 279174
rect 277866 278938 278102 279174
rect 277546 278618 277782 278854
rect 277866 278618 278102 278854
rect 277546 244938 277782 245174
rect 277866 244938 278102 245174
rect 277546 244618 277782 244854
rect 277866 244618 278102 244854
rect 281266 706522 281502 706758
rect 281586 706522 281822 706758
rect 281266 706202 281502 706438
rect 281586 706202 281822 706438
rect 281266 690658 281502 690894
rect 281586 690658 281822 690894
rect 281266 690338 281502 690574
rect 281586 690338 281822 690574
rect 281266 656658 281502 656894
rect 281586 656658 281822 656894
rect 281266 656338 281502 656574
rect 281586 656338 281822 656574
rect 281266 622658 281502 622894
rect 281586 622658 281822 622894
rect 281266 622338 281502 622574
rect 281586 622338 281822 622574
rect 281266 588658 281502 588894
rect 281586 588658 281822 588894
rect 281266 588338 281502 588574
rect 281586 588338 281822 588574
rect 281266 554658 281502 554894
rect 281586 554658 281822 554894
rect 281266 554338 281502 554574
rect 281586 554338 281822 554574
rect 281266 520658 281502 520894
rect 281586 520658 281822 520894
rect 281266 520338 281502 520574
rect 281586 520338 281822 520574
rect 281266 486658 281502 486894
rect 281586 486658 281822 486894
rect 281266 486338 281502 486574
rect 281586 486338 281822 486574
rect 281266 452658 281502 452894
rect 281586 452658 281822 452894
rect 281266 452338 281502 452574
rect 281586 452338 281822 452574
rect 281266 418658 281502 418894
rect 281586 418658 281822 418894
rect 281266 418338 281502 418574
rect 281586 418338 281822 418574
rect 281266 384658 281502 384894
rect 281586 384658 281822 384894
rect 281266 384338 281502 384574
rect 281586 384338 281822 384574
rect 281266 350658 281502 350894
rect 281586 350658 281822 350894
rect 281266 350338 281502 350574
rect 281586 350338 281822 350574
rect 281266 316658 281502 316894
rect 281586 316658 281822 316894
rect 281266 316338 281502 316574
rect 281586 316338 281822 316574
rect 281266 282658 281502 282894
rect 281586 282658 281822 282894
rect 281266 282338 281502 282574
rect 281586 282338 281822 282574
rect 281266 248658 281502 248894
rect 281586 248658 281822 248894
rect 281266 248338 281502 248574
rect 281586 248338 281822 248574
rect 250986 218378 251222 218614
rect 251306 218378 251542 218614
rect 250986 218058 251222 218294
rect 251306 218058 251542 218294
rect 220706 188098 220942 188334
rect 221026 188098 221262 188334
rect 220706 187778 220942 188014
rect 221026 187778 221262 188014
rect 220706 154098 220942 154334
rect 221026 154098 221262 154334
rect 220706 153778 220942 154014
rect 221026 153778 221262 154014
rect 220706 120098 220942 120334
rect 221026 120098 221262 120334
rect 220706 119778 220942 120014
rect 221026 119778 221262 120014
rect 220706 86098 220942 86334
rect 221026 86098 221262 86334
rect 220706 85778 220942 86014
rect 221026 85778 221262 86014
rect 220706 52098 220942 52334
rect 221026 52098 221262 52334
rect 220706 51778 220942 52014
rect 221026 51778 221262 52014
rect 220706 18098 220942 18334
rect 221026 18098 221262 18334
rect 220706 17778 220942 18014
rect 221026 17778 221262 18014
rect 220706 -4422 220942 -4186
rect 221026 -4422 221262 -4186
rect 220706 -4742 220942 -4506
rect 221026 -4742 221262 -4506
rect 224426 191818 224662 192054
rect 224746 191818 224982 192054
rect 224426 191498 224662 191734
rect 224746 191498 224982 191734
rect 224426 157818 224662 158054
rect 224746 157818 224982 158054
rect 224426 157498 224662 157734
rect 224746 157498 224982 157734
rect 224426 123818 224662 124054
rect 224746 123818 224982 124054
rect 224426 123498 224662 123734
rect 224746 123498 224982 123734
rect 224426 89818 224662 90054
rect 224746 89818 224982 90054
rect 224426 89498 224662 89734
rect 224746 89498 224982 89734
rect 224426 55818 224662 56054
rect 224746 55818 224982 56054
rect 224426 55498 224662 55734
rect 224746 55498 224982 55734
rect 224426 21818 224662 22054
rect 224746 21818 224982 22054
rect 224426 21498 224662 21734
rect 224746 21498 224982 21734
rect 224426 -5382 224662 -5146
rect 224746 -5382 224982 -5146
rect 224426 -5702 224662 -5466
rect 224746 -5702 224982 -5466
rect 228146 195538 228382 195774
rect 228466 195538 228702 195774
rect 228146 195218 228382 195454
rect 228466 195218 228702 195454
rect 228146 161538 228382 161774
rect 228466 161538 228702 161774
rect 228146 161218 228382 161454
rect 228466 161218 228702 161454
rect 228146 127538 228382 127774
rect 228466 127538 228702 127774
rect 228146 127218 228382 127454
rect 228466 127218 228702 127454
rect 228146 93538 228382 93774
rect 228466 93538 228702 93774
rect 228146 93218 228382 93454
rect 228466 93218 228702 93454
rect 228146 59538 228382 59774
rect 228466 59538 228702 59774
rect 228146 59218 228382 59454
rect 228466 59218 228702 59454
rect 228146 25538 228382 25774
rect 228466 25538 228702 25774
rect 228146 25218 228382 25454
rect 228466 25218 228702 25454
rect 228146 -6342 228382 -6106
rect 228466 -6342 228702 -6106
rect 228146 -6662 228382 -6426
rect 228466 -6662 228702 -6426
rect 231866 199258 232102 199494
rect 232186 199258 232422 199494
rect 231866 198938 232102 199174
rect 232186 198938 232422 199174
rect 231866 165258 232102 165494
rect 232186 165258 232422 165494
rect 231866 164938 232102 165174
rect 232186 164938 232422 165174
rect 231866 131258 232102 131494
rect 232186 131258 232422 131494
rect 231866 130938 232102 131174
rect 232186 130938 232422 131174
rect 231866 97258 232102 97494
rect 232186 97258 232422 97494
rect 231866 96938 232102 97174
rect 232186 96938 232422 97174
rect 231866 63258 232102 63494
rect 232186 63258 232422 63494
rect 231866 62938 232102 63174
rect 232186 62938 232422 63174
rect 231866 29258 232102 29494
rect 232186 29258 232422 29494
rect 231866 28938 232102 29174
rect 232186 28938 232422 29174
rect 231866 -7302 232102 -7066
rect 232186 -7302 232422 -7066
rect 231866 -7622 232102 -7386
rect 232186 -7622 232422 -7386
rect 239826 207218 240062 207454
rect 240146 207218 240382 207454
rect 239826 206898 240062 207134
rect 240146 206898 240382 207134
rect 239826 173218 240062 173454
rect 240146 173218 240382 173454
rect 239826 172898 240062 173134
rect 240146 172898 240382 173134
rect 239826 139218 240062 139454
rect 240146 139218 240382 139454
rect 239826 138898 240062 139134
rect 240146 138898 240382 139134
rect 239826 105218 240062 105454
rect 240146 105218 240382 105454
rect 239826 104898 240062 105134
rect 240146 104898 240382 105134
rect 239826 71218 240062 71454
rect 240146 71218 240382 71454
rect 239826 70898 240062 71134
rect 240146 70898 240382 71134
rect 239826 37218 240062 37454
rect 240146 37218 240382 37454
rect 239826 36898 240062 37134
rect 240146 36898 240382 37134
rect 239826 3218 240062 3454
rect 240146 3218 240382 3454
rect 239826 2898 240062 3134
rect 240146 2898 240382 3134
rect 239826 -582 240062 -346
rect 240146 -582 240382 -346
rect 239826 -902 240062 -666
rect 240146 -902 240382 -666
rect 243546 210938 243782 211174
rect 243866 210938 244102 211174
rect 243546 210618 243782 210854
rect 243866 210618 244102 210854
rect 243546 176938 243782 177174
rect 243866 176938 244102 177174
rect 243546 176618 243782 176854
rect 243866 176618 244102 176854
rect 243546 142938 243782 143174
rect 243866 142938 244102 143174
rect 243546 142618 243782 142854
rect 243866 142618 244102 142854
rect 243546 108938 243782 109174
rect 243866 108938 244102 109174
rect 243546 108618 243782 108854
rect 243866 108618 244102 108854
rect 243546 74938 243782 75174
rect 243866 74938 244102 75174
rect 243546 74618 243782 74854
rect 243866 74618 244102 74854
rect 243546 40938 243782 41174
rect 243866 40938 244102 41174
rect 243546 40618 243782 40854
rect 243866 40618 244102 40854
rect 243546 6938 243782 7174
rect 243866 6938 244102 7174
rect 243546 6618 243782 6854
rect 243866 6618 244102 6854
rect 243546 -1542 243782 -1306
rect 243866 -1542 244102 -1306
rect 243546 -1862 243782 -1626
rect 243866 -1862 244102 -1626
rect 247266 180658 247502 180894
rect 247586 180658 247822 180894
rect 247266 180338 247502 180574
rect 247586 180338 247822 180574
rect 247266 146658 247502 146894
rect 247586 146658 247822 146894
rect 247266 146338 247502 146574
rect 247586 146338 247822 146574
rect 247266 112658 247502 112894
rect 247586 112658 247822 112894
rect 247266 112338 247502 112574
rect 247586 112338 247822 112574
rect 247266 78658 247502 78894
rect 247586 78658 247822 78894
rect 247266 78338 247502 78574
rect 247586 78338 247822 78574
rect 247266 44658 247502 44894
rect 247586 44658 247822 44894
rect 247266 44338 247502 44574
rect 247586 44338 247822 44574
rect 247266 10658 247502 10894
rect 247586 10658 247822 10894
rect 247266 10338 247502 10574
rect 247586 10338 247822 10574
rect 247266 -2502 247502 -2266
rect 247586 -2502 247822 -2266
rect 247266 -2822 247502 -2586
rect 247586 -2822 247822 -2586
rect 284986 707482 285222 707718
rect 285306 707482 285542 707718
rect 284986 707162 285222 707398
rect 285306 707162 285542 707398
rect 284986 694378 285222 694614
rect 285306 694378 285542 694614
rect 284986 694058 285222 694294
rect 285306 694058 285542 694294
rect 284986 660378 285222 660614
rect 285306 660378 285542 660614
rect 284986 660058 285222 660294
rect 285306 660058 285542 660294
rect 284986 626378 285222 626614
rect 285306 626378 285542 626614
rect 284986 626058 285222 626294
rect 285306 626058 285542 626294
rect 284986 592378 285222 592614
rect 285306 592378 285542 592614
rect 284986 592058 285222 592294
rect 285306 592058 285542 592294
rect 284986 558378 285222 558614
rect 285306 558378 285542 558614
rect 284986 558058 285222 558294
rect 285306 558058 285542 558294
rect 284986 524378 285222 524614
rect 285306 524378 285542 524614
rect 284986 524058 285222 524294
rect 285306 524058 285542 524294
rect 284986 490378 285222 490614
rect 285306 490378 285542 490614
rect 284986 490058 285222 490294
rect 285306 490058 285542 490294
rect 284986 456378 285222 456614
rect 285306 456378 285542 456614
rect 284986 456058 285222 456294
rect 285306 456058 285542 456294
rect 284986 422378 285222 422614
rect 285306 422378 285542 422614
rect 284986 422058 285222 422294
rect 285306 422058 285542 422294
rect 284986 388378 285222 388614
rect 285306 388378 285542 388614
rect 284986 388058 285222 388294
rect 285306 388058 285542 388294
rect 284986 354378 285222 354614
rect 285306 354378 285542 354614
rect 284986 354058 285222 354294
rect 285306 354058 285542 354294
rect 284986 320378 285222 320614
rect 285306 320378 285542 320614
rect 284986 320058 285222 320294
rect 285306 320058 285542 320294
rect 284986 286378 285222 286614
rect 285306 286378 285542 286614
rect 284986 286058 285222 286294
rect 285306 286058 285542 286294
rect 284986 252378 285222 252614
rect 285306 252378 285542 252614
rect 284986 252058 285222 252294
rect 285306 252058 285542 252294
rect 288706 708442 288942 708678
rect 289026 708442 289262 708678
rect 288706 708122 288942 708358
rect 289026 708122 289262 708358
rect 288706 698098 288942 698334
rect 289026 698098 289262 698334
rect 288706 697778 288942 698014
rect 289026 697778 289262 698014
rect 288706 664098 288942 664334
rect 289026 664098 289262 664334
rect 288706 663778 288942 664014
rect 289026 663778 289262 664014
rect 288706 630098 288942 630334
rect 289026 630098 289262 630334
rect 288706 629778 288942 630014
rect 289026 629778 289262 630014
rect 288706 596098 288942 596334
rect 289026 596098 289262 596334
rect 288706 595778 288942 596014
rect 289026 595778 289262 596014
rect 288706 562098 288942 562334
rect 289026 562098 289262 562334
rect 288706 561778 288942 562014
rect 289026 561778 289262 562014
rect 288706 528098 288942 528334
rect 289026 528098 289262 528334
rect 288706 527778 288942 528014
rect 289026 527778 289262 528014
rect 288706 494098 288942 494334
rect 289026 494098 289262 494334
rect 288706 493778 288942 494014
rect 289026 493778 289262 494014
rect 288706 460098 288942 460334
rect 289026 460098 289262 460334
rect 288706 459778 288942 460014
rect 289026 459778 289262 460014
rect 288706 426098 288942 426334
rect 289026 426098 289262 426334
rect 288706 425778 288942 426014
rect 289026 425778 289262 426014
rect 288706 392098 288942 392334
rect 289026 392098 289262 392334
rect 288706 391778 288942 392014
rect 289026 391778 289262 392014
rect 288706 358098 288942 358334
rect 289026 358098 289262 358334
rect 288706 357778 288942 358014
rect 289026 357778 289262 358014
rect 288706 324098 288942 324334
rect 289026 324098 289262 324334
rect 288706 323778 288942 324014
rect 289026 323778 289262 324014
rect 288706 290098 288942 290334
rect 289026 290098 289262 290334
rect 288706 289778 288942 290014
rect 289026 289778 289262 290014
rect 288706 256098 288942 256334
rect 289026 256098 289262 256334
rect 288706 255778 288942 256014
rect 289026 255778 289262 256014
rect 292426 709402 292662 709638
rect 292746 709402 292982 709638
rect 292426 709082 292662 709318
rect 292746 709082 292982 709318
rect 292426 667818 292662 668054
rect 292746 667818 292982 668054
rect 292426 667498 292662 667734
rect 292746 667498 292982 667734
rect 292426 633818 292662 634054
rect 292746 633818 292982 634054
rect 292426 633498 292662 633734
rect 292746 633498 292982 633734
rect 292426 599818 292662 600054
rect 292746 599818 292982 600054
rect 292426 599498 292662 599734
rect 292746 599498 292982 599734
rect 292426 565818 292662 566054
rect 292746 565818 292982 566054
rect 292426 565498 292662 565734
rect 292746 565498 292982 565734
rect 292426 531818 292662 532054
rect 292746 531818 292982 532054
rect 292426 531498 292662 531734
rect 292746 531498 292982 531734
rect 292426 497818 292662 498054
rect 292746 497818 292982 498054
rect 292426 497498 292662 497734
rect 292746 497498 292982 497734
rect 292426 463818 292662 464054
rect 292746 463818 292982 464054
rect 292426 463498 292662 463734
rect 292746 463498 292982 463734
rect 292426 429818 292662 430054
rect 292746 429818 292982 430054
rect 292426 429498 292662 429734
rect 292746 429498 292982 429734
rect 292426 395818 292662 396054
rect 292746 395818 292982 396054
rect 292426 395498 292662 395734
rect 292746 395498 292982 395734
rect 292426 361818 292662 362054
rect 292746 361818 292982 362054
rect 292426 361498 292662 361734
rect 292746 361498 292982 361734
rect 292426 327818 292662 328054
rect 292746 327818 292982 328054
rect 292426 327498 292662 327734
rect 292746 327498 292982 327734
rect 292426 293818 292662 294054
rect 292746 293818 292982 294054
rect 292426 293498 292662 293734
rect 292746 293498 292982 293734
rect 292426 259818 292662 260054
rect 292746 259818 292982 260054
rect 292426 259498 292662 259734
rect 292746 259498 292982 259734
rect 292426 225755 292662 225991
rect 292746 225755 292982 225991
rect 296146 710362 296382 710598
rect 296466 710362 296702 710598
rect 296146 710042 296382 710278
rect 296466 710042 296702 710278
rect 296146 671538 296382 671774
rect 296466 671538 296702 671774
rect 296146 671218 296382 671454
rect 296466 671218 296702 671454
rect 296146 637538 296382 637774
rect 296466 637538 296702 637774
rect 296146 637218 296382 637454
rect 296466 637218 296702 637454
rect 296146 603538 296382 603774
rect 296466 603538 296702 603774
rect 296146 603218 296382 603454
rect 296466 603218 296702 603454
rect 296146 569538 296382 569774
rect 296466 569538 296702 569774
rect 296146 569218 296382 569454
rect 296466 569218 296702 569454
rect 296146 535538 296382 535774
rect 296466 535538 296702 535774
rect 296146 535218 296382 535454
rect 296466 535218 296702 535454
rect 296146 501538 296382 501774
rect 296466 501538 296702 501774
rect 296146 501218 296382 501454
rect 296466 501218 296702 501454
rect 296146 467538 296382 467774
rect 296466 467538 296702 467774
rect 296146 467218 296382 467454
rect 296466 467218 296702 467454
rect 296146 433538 296382 433774
rect 296466 433538 296702 433774
rect 296146 433218 296382 433454
rect 296466 433218 296702 433454
rect 296146 399538 296382 399774
rect 296466 399538 296702 399774
rect 296146 399218 296382 399454
rect 296466 399218 296702 399454
rect 296146 365538 296382 365774
rect 296466 365538 296702 365774
rect 296146 365218 296382 365454
rect 296466 365218 296702 365454
rect 296146 331538 296382 331774
rect 296466 331538 296702 331774
rect 296146 331218 296382 331454
rect 296466 331218 296702 331454
rect 296146 297538 296382 297774
rect 296466 297538 296702 297774
rect 296146 297218 296382 297454
rect 296466 297218 296702 297454
rect 296146 263538 296382 263774
rect 296466 263538 296702 263774
rect 296146 263218 296382 263454
rect 296466 263218 296702 263454
rect 296146 229538 296382 229774
rect 296466 229538 296702 229774
rect 296146 229218 296382 229454
rect 296466 229218 296702 229454
rect 299866 711322 300102 711558
rect 300186 711322 300422 711558
rect 299866 711002 300102 711238
rect 300186 711002 300422 711238
rect 299866 675258 300102 675494
rect 300186 675258 300422 675494
rect 299866 674938 300102 675174
rect 300186 674938 300422 675174
rect 299866 641258 300102 641494
rect 300186 641258 300422 641494
rect 299866 640938 300102 641174
rect 300186 640938 300422 641174
rect 299866 607258 300102 607494
rect 300186 607258 300422 607494
rect 299866 606938 300102 607174
rect 300186 606938 300422 607174
rect 299866 573258 300102 573494
rect 300186 573258 300422 573494
rect 299866 572938 300102 573174
rect 300186 572938 300422 573174
rect 299866 539258 300102 539494
rect 300186 539258 300422 539494
rect 299866 538938 300102 539174
rect 300186 538938 300422 539174
rect 299866 505258 300102 505494
rect 300186 505258 300422 505494
rect 299866 504938 300102 505174
rect 300186 504938 300422 505174
rect 299866 471258 300102 471494
rect 300186 471258 300422 471494
rect 299866 470938 300102 471174
rect 300186 470938 300422 471174
rect 299866 437258 300102 437494
rect 300186 437258 300422 437494
rect 299866 436938 300102 437174
rect 300186 436938 300422 437174
rect 299866 403258 300102 403494
rect 300186 403258 300422 403494
rect 299866 402938 300102 403174
rect 300186 402938 300422 403174
rect 299866 369258 300102 369494
rect 300186 369258 300422 369494
rect 299866 368938 300102 369174
rect 300186 368938 300422 369174
rect 299866 335258 300102 335494
rect 300186 335258 300422 335494
rect 299866 334938 300102 335174
rect 300186 334938 300422 335174
rect 299866 301258 300102 301494
rect 300186 301258 300422 301494
rect 299866 300938 300102 301174
rect 300186 300938 300422 301174
rect 299866 267258 300102 267494
rect 300186 267258 300422 267494
rect 299866 266938 300102 267174
rect 300186 266938 300422 267174
rect 299866 233258 300102 233494
rect 300186 233258 300422 233494
rect 299866 232938 300102 233174
rect 300186 232938 300422 233174
rect 307826 704602 308062 704838
rect 308146 704602 308382 704838
rect 307826 704282 308062 704518
rect 308146 704282 308382 704518
rect 307826 683218 308062 683454
rect 308146 683218 308382 683454
rect 307826 682898 308062 683134
rect 308146 682898 308382 683134
rect 307826 649218 308062 649454
rect 308146 649218 308382 649454
rect 307826 648898 308062 649134
rect 308146 648898 308382 649134
rect 307826 615218 308062 615454
rect 308146 615218 308382 615454
rect 307826 614898 308062 615134
rect 308146 614898 308382 615134
rect 307826 581218 308062 581454
rect 308146 581218 308382 581454
rect 307826 580898 308062 581134
rect 308146 580898 308382 581134
rect 307826 547218 308062 547454
rect 308146 547218 308382 547454
rect 307826 546898 308062 547134
rect 308146 546898 308382 547134
rect 307826 513218 308062 513454
rect 308146 513218 308382 513454
rect 307826 512898 308062 513134
rect 308146 512898 308382 513134
rect 307826 479218 308062 479454
rect 308146 479218 308382 479454
rect 307826 478898 308062 479134
rect 308146 478898 308382 479134
rect 307826 445218 308062 445454
rect 308146 445218 308382 445454
rect 307826 444898 308062 445134
rect 308146 444898 308382 445134
rect 307826 411218 308062 411454
rect 308146 411218 308382 411454
rect 307826 410898 308062 411134
rect 308146 410898 308382 411134
rect 307826 377218 308062 377454
rect 308146 377218 308382 377454
rect 307826 376898 308062 377134
rect 308146 376898 308382 377134
rect 307826 343218 308062 343454
rect 308146 343218 308382 343454
rect 307826 342898 308062 343134
rect 308146 342898 308382 343134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 275218 308062 275454
rect 308146 275218 308382 275454
rect 307826 274898 308062 275134
rect 308146 274898 308382 275134
rect 307826 241218 308062 241454
rect 308146 241218 308382 241454
rect 307826 240898 308062 241134
rect 308146 240898 308382 241134
rect 311546 705562 311782 705798
rect 311866 705562 312102 705798
rect 311546 705242 311782 705478
rect 311866 705242 312102 705478
rect 311546 686938 311782 687174
rect 311866 686938 312102 687174
rect 311546 686618 311782 686854
rect 311866 686618 312102 686854
rect 311546 652938 311782 653174
rect 311866 652938 312102 653174
rect 311546 652618 311782 652854
rect 311866 652618 312102 652854
rect 311546 618938 311782 619174
rect 311866 618938 312102 619174
rect 311546 618618 311782 618854
rect 311866 618618 312102 618854
rect 311546 584938 311782 585174
rect 311866 584938 312102 585174
rect 311546 584618 311782 584854
rect 311866 584618 312102 584854
rect 311546 550938 311782 551174
rect 311866 550938 312102 551174
rect 311546 550618 311782 550854
rect 311866 550618 312102 550854
rect 311546 516938 311782 517174
rect 311866 516938 312102 517174
rect 311546 516618 311782 516854
rect 311866 516618 312102 516854
rect 311546 482938 311782 483174
rect 311866 482938 312102 483174
rect 311546 482618 311782 482854
rect 311866 482618 312102 482854
rect 311546 448938 311782 449174
rect 311866 448938 312102 449174
rect 311546 448618 311782 448854
rect 311866 448618 312102 448854
rect 311546 414938 311782 415174
rect 311866 414938 312102 415174
rect 311546 414618 311782 414854
rect 311866 414618 312102 414854
rect 311546 380938 311782 381174
rect 311866 380938 312102 381174
rect 311546 380618 311782 380854
rect 311866 380618 312102 380854
rect 311546 346938 311782 347174
rect 311866 346938 312102 347174
rect 311546 346618 311782 346854
rect 311866 346618 312102 346854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 278938 311782 279174
rect 311866 278938 312102 279174
rect 311546 278618 311782 278854
rect 311866 278618 312102 278854
rect 311546 244938 311782 245174
rect 311866 244938 312102 245174
rect 311546 244618 311782 244854
rect 311866 244618 312102 244854
rect 281266 214658 281502 214894
rect 281586 214658 281822 214894
rect 250986 184378 251222 184614
rect 251306 184378 251542 184614
rect 250986 184058 251222 184294
rect 251306 184058 251542 184294
rect 250986 150378 251222 150614
rect 251306 150378 251542 150614
rect 250986 150058 251222 150294
rect 251306 150058 251542 150294
rect 250986 116378 251222 116614
rect 251306 116378 251542 116614
rect 250986 116058 251222 116294
rect 251306 116058 251542 116294
rect 250986 82378 251222 82614
rect 251306 82378 251542 82614
rect 250986 82058 251222 82294
rect 251306 82058 251542 82294
rect 250986 48378 251222 48614
rect 251306 48378 251542 48614
rect 250986 48058 251222 48294
rect 251306 48058 251542 48294
rect 250986 14378 251222 14614
rect 251306 14378 251542 14614
rect 250986 14058 251222 14294
rect 251306 14058 251542 14294
rect 250986 -3462 251222 -3226
rect 251306 -3462 251542 -3226
rect 250986 -3782 251222 -3546
rect 251306 -3782 251542 -3546
rect 254706 188098 254942 188334
rect 255026 188098 255262 188334
rect 254706 187778 254942 188014
rect 255026 187778 255262 188014
rect 254706 154098 254942 154334
rect 255026 154098 255262 154334
rect 254706 153778 254942 154014
rect 255026 153778 255262 154014
rect 254706 120098 254942 120334
rect 255026 120098 255262 120334
rect 254706 119778 254942 120014
rect 255026 119778 255262 120014
rect 254706 86098 254942 86334
rect 255026 86098 255262 86334
rect 254706 85778 254942 86014
rect 255026 85778 255262 86014
rect 254706 52098 254942 52334
rect 255026 52098 255262 52334
rect 254706 51778 254942 52014
rect 255026 51778 255262 52014
rect 254706 18098 254942 18334
rect 255026 18098 255262 18334
rect 254706 17778 254942 18014
rect 255026 17778 255262 18014
rect 254706 -4422 254942 -4186
rect 255026 -4422 255262 -4186
rect 254706 -4742 254942 -4506
rect 255026 -4742 255262 -4506
rect 258426 191818 258662 192054
rect 258746 191818 258982 192054
rect 258426 191498 258662 191734
rect 258746 191498 258982 191734
rect 258426 157818 258662 158054
rect 258746 157818 258982 158054
rect 258426 157498 258662 157734
rect 258746 157498 258982 157734
rect 258426 123818 258662 124054
rect 258746 123818 258982 124054
rect 258426 123498 258662 123734
rect 258746 123498 258982 123734
rect 258426 89818 258662 90054
rect 258746 89818 258982 90054
rect 258426 89498 258662 89734
rect 258746 89498 258982 89734
rect 258426 55818 258662 56054
rect 258746 55818 258982 56054
rect 258426 55498 258662 55734
rect 258746 55498 258982 55734
rect 258426 21818 258662 22054
rect 258746 21818 258982 22054
rect 258426 21498 258662 21734
rect 258746 21498 258982 21734
rect 258426 -5382 258662 -5146
rect 258746 -5382 258982 -5146
rect 258426 -5702 258662 -5466
rect 258746 -5702 258982 -5466
rect 262146 195538 262382 195774
rect 262466 195538 262702 195774
rect 262146 195218 262382 195454
rect 262466 195218 262702 195454
rect 262146 161538 262382 161774
rect 262466 161538 262702 161774
rect 262146 161218 262382 161454
rect 262466 161218 262702 161454
rect 262146 127538 262382 127774
rect 262466 127538 262702 127774
rect 262146 127218 262382 127454
rect 262466 127218 262702 127454
rect 262146 93538 262382 93774
rect 262466 93538 262702 93774
rect 262146 93218 262382 93454
rect 262466 93218 262702 93454
rect 262146 59538 262382 59774
rect 262466 59538 262702 59774
rect 262146 59218 262382 59454
rect 262466 59218 262702 59454
rect 262146 25538 262382 25774
rect 262466 25538 262702 25774
rect 262146 25218 262382 25454
rect 262466 25218 262702 25454
rect 262146 -6342 262382 -6106
rect 262466 -6342 262702 -6106
rect 262146 -6662 262382 -6426
rect 262466 -6662 262702 -6426
rect 265866 199258 266102 199494
rect 266186 199258 266422 199494
rect 265866 198938 266102 199174
rect 266186 198938 266422 199174
rect 265866 165258 266102 165494
rect 266186 165258 266422 165494
rect 265866 164938 266102 165174
rect 266186 164938 266422 165174
rect 265866 131258 266102 131494
rect 266186 131258 266422 131494
rect 265866 130938 266102 131174
rect 266186 130938 266422 131174
rect 265866 97258 266102 97494
rect 266186 97258 266422 97494
rect 265866 96938 266102 97174
rect 266186 96938 266422 97174
rect 265866 63258 266102 63494
rect 266186 63258 266422 63494
rect 265866 62938 266102 63174
rect 266186 62938 266422 63174
rect 265866 29258 266102 29494
rect 266186 29258 266422 29494
rect 265866 28938 266102 29174
rect 266186 28938 266422 29174
rect 265866 -7302 266102 -7066
rect 266186 -7302 266422 -7066
rect 265866 -7622 266102 -7386
rect 266186 -7622 266422 -7386
rect 273826 207218 274062 207454
rect 274146 207218 274382 207454
rect 273826 206898 274062 207134
rect 274146 206898 274382 207134
rect 273826 173218 274062 173454
rect 274146 173218 274382 173454
rect 273826 172898 274062 173134
rect 274146 172898 274382 173134
rect 273826 139218 274062 139454
rect 274146 139218 274382 139454
rect 273826 138898 274062 139134
rect 274146 138898 274382 139134
rect 273826 105218 274062 105454
rect 274146 105218 274382 105454
rect 273826 104898 274062 105134
rect 274146 104898 274382 105134
rect 273826 71218 274062 71454
rect 274146 71218 274382 71454
rect 273826 70898 274062 71134
rect 274146 70898 274382 71134
rect 273826 37218 274062 37454
rect 274146 37218 274382 37454
rect 273826 36898 274062 37134
rect 274146 36898 274382 37134
rect 273826 3218 274062 3454
rect 274146 3218 274382 3454
rect 273826 2898 274062 3134
rect 274146 2898 274382 3134
rect 273826 -582 274062 -346
rect 274146 -582 274382 -346
rect 273826 -902 274062 -666
rect 274146 -902 274382 -666
rect 277546 210938 277782 211174
rect 277866 210938 278102 211174
rect 277546 210618 277782 210854
rect 277866 210618 278102 210854
rect 277546 176938 277782 177174
rect 277866 176938 278102 177174
rect 277546 176618 277782 176854
rect 277866 176618 278102 176854
rect 277546 142938 277782 143174
rect 277866 142938 278102 143174
rect 277546 142618 277782 142854
rect 277866 142618 278102 142854
rect 277546 108938 277782 109174
rect 277866 108938 278102 109174
rect 277546 108618 277782 108854
rect 277866 108618 278102 108854
rect 277546 74938 277782 75174
rect 277866 74938 278102 75174
rect 277546 74618 277782 74854
rect 277866 74618 278102 74854
rect 277546 40938 277782 41174
rect 277866 40938 278102 41174
rect 277546 40618 277782 40854
rect 277866 40618 278102 40854
rect 277546 6938 277782 7174
rect 277866 6938 278102 7174
rect 277546 6618 277782 6854
rect 277866 6618 278102 6854
rect 277546 -1542 277782 -1306
rect 277866 -1542 278102 -1306
rect 277546 -1862 277782 -1626
rect 277866 -1862 278102 -1626
rect 281266 214338 281502 214574
rect 281586 214338 281822 214574
rect 281266 180658 281502 180894
rect 281586 180658 281822 180894
rect 281266 180338 281502 180574
rect 281586 180338 281822 180574
rect 281266 146658 281502 146894
rect 281586 146658 281822 146894
rect 281266 146338 281502 146574
rect 281586 146338 281822 146574
rect 281266 112658 281502 112894
rect 281586 112658 281822 112894
rect 281266 112338 281502 112574
rect 281586 112338 281822 112574
rect 281266 78658 281502 78894
rect 281586 78658 281822 78894
rect 281266 78338 281502 78574
rect 281586 78338 281822 78574
rect 281266 44658 281502 44894
rect 281586 44658 281822 44894
rect 281266 44338 281502 44574
rect 281586 44338 281822 44574
rect 281266 10658 281502 10894
rect 281586 10658 281822 10894
rect 281266 10338 281502 10574
rect 281586 10338 281822 10574
rect 281266 -2502 281502 -2266
rect 281586 -2502 281822 -2266
rect 281266 -2822 281502 -2586
rect 281586 -2822 281822 -2586
rect 284986 184378 285222 184614
rect 285306 184378 285542 184614
rect 284986 184058 285222 184294
rect 285306 184058 285542 184294
rect 284986 150378 285222 150614
rect 285306 150378 285542 150614
rect 284986 150058 285222 150294
rect 285306 150058 285542 150294
rect 284986 116378 285222 116614
rect 285306 116378 285542 116614
rect 284986 116058 285222 116294
rect 285306 116058 285542 116294
rect 284986 82378 285222 82614
rect 285306 82378 285542 82614
rect 284986 82058 285222 82294
rect 285306 82058 285542 82294
rect 284986 48378 285222 48614
rect 285306 48378 285542 48614
rect 284986 48058 285222 48294
rect 285306 48058 285542 48294
rect 284986 14378 285222 14614
rect 285306 14378 285542 14614
rect 284986 14058 285222 14294
rect 285306 14058 285542 14294
rect 284986 -3462 285222 -3226
rect 285306 -3462 285542 -3226
rect 284986 -3782 285222 -3546
rect 285306 -3782 285542 -3546
rect 288706 188098 288942 188334
rect 289026 188098 289262 188334
rect 288706 187778 288942 188014
rect 289026 187778 289262 188014
rect 288706 154098 288942 154334
rect 289026 154098 289262 154334
rect 288706 153778 288942 154014
rect 289026 153778 289262 154014
rect 288706 120098 288942 120334
rect 289026 120098 289262 120334
rect 288706 119778 288942 120014
rect 289026 119778 289262 120014
rect 288706 86098 288942 86334
rect 289026 86098 289262 86334
rect 288706 85778 288942 86014
rect 289026 85778 289262 86014
rect 288706 52098 288942 52334
rect 289026 52098 289262 52334
rect 288706 51778 288942 52014
rect 289026 51778 289262 52014
rect 288706 18098 288942 18334
rect 289026 18098 289262 18334
rect 288706 17778 288942 18014
rect 289026 17778 289262 18014
rect 288706 -4422 288942 -4186
rect 289026 -4422 289262 -4186
rect 288706 -4742 288942 -4506
rect 289026 -4742 289262 -4506
rect 292426 191818 292662 192054
rect 292746 191818 292982 192054
rect 292426 191498 292662 191734
rect 292746 191498 292982 191734
rect 292426 157818 292662 158054
rect 292746 157818 292982 158054
rect 292426 157498 292662 157734
rect 292746 157498 292982 157734
rect 292426 123818 292662 124054
rect 292746 123818 292982 124054
rect 292426 123498 292662 123734
rect 292746 123498 292982 123734
rect 292426 89818 292662 90054
rect 292746 89818 292982 90054
rect 292426 89498 292662 89734
rect 292746 89498 292982 89734
rect 292426 55818 292662 56054
rect 292746 55818 292982 56054
rect 292426 55498 292662 55734
rect 292746 55498 292982 55734
rect 292426 21818 292662 22054
rect 292746 21818 292982 22054
rect 292426 21498 292662 21734
rect 292746 21498 292982 21734
rect 292426 -5382 292662 -5146
rect 292746 -5382 292982 -5146
rect 292426 -5702 292662 -5466
rect 292746 -5702 292982 -5466
rect 296146 195538 296382 195774
rect 296466 195538 296702 195774
rect 296146 195218 296382 195454
rect 296466 195218 296702 195454
rect 296146 161538 296382 161774
rect 296466 161538 296702 161774
rect 296146 161218 296382 161454
rect 296466 161218 296702 161454
rect 296146 127538 296382 127774
rect 296466 127538 296702 127774
rect 296146 127218 296382 127454
rect 296466 127218 296702 127454
rect 296146 93538 296382 93774
rect 296466 93538 296702 93774
rect 296146 93218 296382 93454
rect 296466 93218 296702 93454
rect 296146 59538 296382 59774
rect 296466 59538 296702 59774
rect 296146 59218 296382 59454
rect 296466 59218 296702 59454
rect 296146 25538 296382 25774
rect 296466 25538 296702 25774
rect 296146 25218 296382 25454
rect 296466 25218 296702 25454
rect 296146 -6342 296382 -6106
rect 296466 -6342 296702 -6106
rect 296146 -6662 296382 -6426
rect 296466 -6662 296702 -6426
rect 299866 199258 300102 199494
rect 300186 199258 300422 199494
rect 299866 198938 300102 199174
rect 300186 198938 300422 199174
rect 299866 165258 300102 165494
rect 300186 165258 300422 165494
rect 299866 164938 300102 165174
rect 300186 164938 300422 165174
rect 299866 131258 300102 131494
rect 300186 131258 300422 131494
rect 299866 130938 300102 131174
rect 300186 130938 300422 131174
rect 299866 97258 300102 97494
rect 300186 97258 300422 97494
rect 299866 96938 300102 97174
rect 300186 96938 300422 97174
rect 299866 63258 300102 63494
rect 300186 63258 300422 63494
rect 299866 62938 300102 63174
rect 300186 62938 300422 63174
rect 299866 29258 300102 29494
rect 300186 29258 300422 29494
rect 299866 28938 300102 29174
rect 300186 28938 300422 29174
rect 299866 -7302 300102 -7066
rect 300186 -7302 300422 -7066
rect 299866 -7622 300102 -7386
rect 300186 -7622 300422 -7386
rect 307826 207218 308062 207454
rect 308146 207218 308382 207454
rect 307826 206898 308062 207134
rect 308146 206898 308382 207134
rect 307826 173218 308062 173454
rect 308146 173218 308382 173454
rect 307826 172898 308062 173134
rect 308146 172898 308382 173134
rect 307826 139218 308062 139454
rect 308146 139218 308382 139454
rect 307826 138898 308062 139134
rect 308146 138898 308382 139134
rect 307826 105218 308062 105454
rect 308146 105218 308382 105454
rect 307826 104898 308062 105134
rect 308146 104898 308382 105134
rect 307826 71218 308062 71454
rect 308146 71218 308382 71454
rect 307826 70898 308062 71134
rect 308146 70898 308382 71134
rect 307826 37218 308062 37454
rect 308146 37218 308382 37454
rect 307826 36898 308062 37134
rect 308146 36898 308382 37134
rect 307826 3218 308062 3454
rect 308146 3218 308382 3454
rect 307826 2898 308062 3134
rect 308146 2898 308382 3134
rect 307826 -582 308062 -346
rect 308146 -582 308382 -346
rect 307826 -902 308062 -666
rect 308146 -902 308382 -666
rect 315266 706522 315502 706758
rect 315586 706522 315822 706758
rect 315266 706202 315502 706438
rect 315586 706202 315822 706438
rect 315266 690658 315502 690894
rect 315586 690658 315822 690894
rect 315266 690338 315502 690574
rect 315586 690338 315822 690574
rect 315266 656658 315502 656894
rect 315586 656658 315822 656894
rect 315266 656338 315502 656574
rect 315586 656338 315822 656574
rect 315266 622658 315502 622894
rect 315586 622658 315822 622894
rect 315266 622338 315502 622574
rect 315586 622338 315822 622574
rect 315266 588658 315502 588894
rect 315586 588658 315822 588894
rect 315266 588338 315502 588574
rect 315586 588338 315822 588574
rect 315266 554658 315502 554894
rect 315586 554658 315822 554894
rect 315266 554338 315502 554574
rect 315586 554338 315822 554574
rect 315266 520658 315502 520894
rect 315586 520658 315822 520894
rect 315266 520338 315502 520574
rect 315586 520338 315822 520574
rect 315266 486658 315502 486894
rect 315586 486658 315822 486894
rect 315266 486338 315502 486574
rect 315586 486338 315822 486574
rect 315266 452658 315502 452894
rect 315586 452658 315822 452894
rect 315266 452338 315502 452574
rect 315586 452338 315822 452574
rect 315266 418658 315502 418894
rect 315586 418658 315822 418894
rect 315266 418338 315502 418574
rect 315586 418338 315822 418574
rect 315266 384658 315502 384894
rect 315586 384658 315822 384894
rect 315266 384338 315502 384574
rect 315586 384338 315822 384574
rect 315266 350658 315502 350894
rect 315586 350658 315822 350894
rect 315266 350338 315502 350574
rect 315586 350338 315822 350574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 282658 315502 282894
rect 315586 282658 315822 282894
rect 315266 282338 315502 282574
rect 315586 282338 315822 282574
rect 315266 248658 315502 248894
rect 315586 248658 315822 248894
rect 315266 248338 315502 248574
rect 315586 248338 315822 248574
rect 318986 707482 319222 707718
rect 319306 707482 319542 707718
rect 318986 707162 319222 707398
rect 319306 707162 319542 707398
rect 318986 694378 319222 694614
rect 319306 694378 319542 694614
rect 318986 694058 319222 694294
rect 319306 694058 319542 694294
rect 318986 660378 319222 660614
rect 319306 660378 319542 660614
rect 318986 660058 319222 660294
rect 319306 660058 319542 660294
rect 318986 626378 319222 626614
rect 319306 626378 319542 626614
rect 318986 626058 319222 626294
rect 319306 626058 319542 626294
rect 318986 592378 319222 592614
rect 319306 592378 319542 592614
rect 318986 592058 319222 592294
rect 319306 592058 319542 592294
rect 318986 558378 319222 558614
rect 319306 558378 319542 558614
rect 318986 558058 319222 558294
rect 319306 558058 319542 558294
rect 318986 524378 319222 524614
rect 319306 524378 319542 524614
rect 318986 524058 319222 524294
rect 319306 524058 319542 524294
rect 318986 490378 319222 490614
rect 319306 490378 319542 490614
rect 318986 490058 319222 490294
rect 319306 490058 319542 490294
rect 318986 456378 319222 456614
rect 319306 456378 319542 456614
rect 318986 456058 319222 456294
rect 319306 456058 319542 456294
rect 318986 422378 319222 422614
rect 319306 422378 319542 422614
rect 318986 422058 319222 422294
rect 319306 422058 319542 422294
rect 318986 388378 319222 388614
rect 319306 388378 319542 388614
rect 318986 388058 319222 388294
rect 319306 388058 319542 388294
rect 318986 354378 319222 354614
rect 319306 354378 319542 354614
rect 318986 354058 319222 354294
rect 319306 354058 319542 354294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 286378 319222 286614
rect 319306 286378 319542 286614
rect 318986 286058 319222 286294
rect 319306 286058 319542 286294
rect 318986 252378 319222 252614
rect 319306 252378 319542 252614
rect 318986 252058 319222 252294
rect 319306 252058 319542 252294
rect 322706 708442 322942 708678
rect 323026 708442 323262 708678
rect 322706 708122 322942 708358
rect 323026 708122 323262 708358
rect 322706 698098 322942 698334
rect 323026 698098 323262 698334
rect 322706 697778 322942 698014
rect 323026 697778 323262 698014
rect 322706 664098 322942 664334
rect 323026 664098 323262 664334
rect 322706 663778 322942 664014
rect 323026 663778 323262 664014
rect 322706 630098 322942 630334
rect 323026 630098 323262 630334
rect 322706 629778 322942 630014
rect 323026 629778 323262 630014
rect 322706 596098 322942 596334
rect 323026 596098 323262 596334
rect 322706 595778 322942 596014
rect 323026 595778 323262 596014
rect 322706 562098 322942 562334
rect 323026 562098 323262 562334
rect 322706 561778 322942 562014
rect 323026 561778 323262 562014
rect 322706 528098 322942 528334
rect 323026 528098 323262 528334
rect 322706 527778 322942 528014
rect 323026 527778 323262 528014
rect 322706 494098 322942 494334
rect 323026 494098 323262 494334
rect 322706 493778 322942 494014
rect 323026 493778 323262 494014
rect 322706 460098 322942 460334
rect 323026 460098 323262 460334
rect 322706 459778 322942 460014
rect 323026 459778 323262 460014
rect 322706 426098 322942 426334
rect 323026 426098 323262 426334
rect 322706 425778 322942 426014
rect 323026 425778 323262 426014
rect 322706 392098 322942 392334
rect 323026 392098 323262 392334
rect 322706 391778 322942 392014
rect 323026 391778 323262 392014
rect 322706 358098 322942 358334
rect 323026 358098 323262 358334
rect 322706 357778 322942 358014
rect 323026 357778 323262 358014
rect 322706 324098 322942 324334
rect 323026 324098 323262 324334
rect 322706 323778 322942 324014
rect 323026 323778 323262 324014
rect 322706 290098 322942 290334
rect 323026 290098 323262 290334
rect 322706 289778 322942 290014
rect 323026 289778 323262 290014
rect 322706 256098 322942 256334
rect 323026 256098 323262 256334
rect 322706 255778 322942 256014
rect 323026 255778 323262 256014
rect 326426 709402 326662 709638
rect 326746 709402 326982 709638
rect 326426 709082 326662 709318
rect 326746 709082 326982 709318
rect 326426 667818 326662 668054
rect 326746 667818 326982 668054
rect 326426 667498 326662 667734
rect 326746 667498 326982 667734
rect 326426 633818 326662 634054
rect 326746 633818 326982 634054
rect 326426 633498 326662 633734
rect 326746 633498 326982 633734
rect 326426 599818 326662 600054
rect 326746 599818 326982 600054
rect 326426 599498 326662 599734
rect 326746 599498 326982 599734
rect 326426 565818 326662 566054
rect 326746 565818 326982 566054
rect 326426 565498 326662 565734
rect 326746 565498 326982 565734
rect 326426 531818 326662 532054
rect 326746 531818 326982 532054
rect 326426 531498 326662 531734
rect 326746 531498 326982 531734
rect 326426 497818 326662 498054
rect 326746 497818 326982 498054
rect 326426 497498 326662 497734
rect 326746 497498 326982 497734
rect 326426 463818 326662 464054
rect 326746 463818 326982 464054
rect 326426 463498 326662 463734
rect 326746 463498 326982 463734
rect 326426 429818 326662 430054
rect 326746 429818 326982 430054
rect 326426 429498 326662 429734
rect 326746 429498 326982 429734
rect 326426 395818 326662 396054
rect 326746 395818 326982 396054
rect 326426 395498 326662 395734
rect 326746 395498 326982 395734
rect 326426 361818 326662 362054
rect 326746 361818 326982 362054
rect 326426 361498 326662 361734
rect 326746 361498 326982 361734
rect 326426 327818 326662 328054
rect 326746 327818 326982 328054
rect 326426 327498 326662 327734
rect 326746 327498 326982 327734
rect 326426 293818 326662 294054
rect 326746 293818 326982 294054
rect 326426 293498 326662 293734
rect 326746 293498 326982 293734
rect 326426 259818 326662 260054
rect 326746 259818 326982 260054
rect 326426 259498 326662 259734
rect 326746 259498 326982 259734
rect 326426 225755 326662 225991
rect 326746 225755 326982 225991
rect 330146 710362 330382 710598
rect 330466 710362 330702 710598
rect 330146 710042 330382 710278
rect 330466 710042 330702 710278
rect 330146 671538 330382 671774
rect 330466 671538 330702 671774
rect 330146 671218 330382 671454
rect 330466 671218 330702 671454
rect 330146 637538 330382 637774
rect 330466 637538 330702 637774
rect 330146 637218 330382 637454
rect 330466 637218 330702 637454
rect 330146 603538 330382 603774
rect 330466 603538 330702 603774
rect 330146 603218 330382 603454
rect 330466 603218 330702 603454
rect 330146 569538 330382 569774
rect 330466 569538 330702 569774
rect 330146 569218 330382 569454
rect 330466 569218 330702 569454
rect 330146 535538 330382 535774
rect 330466 535538 330702 535774
rect 330146 535218 330382 535454
rect 330466 535218 330702 535454
rect 330146 501538 330382 501774
rect 330466 501538 330702 501774
rect 330146 501218 330382 501454
rect 330466 501218 330702 501454
rect 330146 467538 330382 467774
rect 330466 467538 330702 467774
rect 330146 467218 330382 467454
rect 330466 467218 330702 467454
rect 330146 433538 330382 433774
rect 330466 433538 330702 433774
rect 330146 433218 330382 433454
rect 330466 433218 330702 433454
rect 330146 399538 330382 399774
rect 330466 399538 330702 399774
rect 330146 399218 330382 399454
rect 330466 399218 330702 399454
rect 330146 365538 330382 365774
rect 330466 365538 330702 365774
rect 330146 365218 330382 365454
rect 330466 365218 330702 365454
rect 330146 331538 330382 331774
rect 330466 331538 330702 331774
rect 330146 331218 330382 331454
rect 330466 331218 330702 331454
rect 330146 297538 330382 297774
rect 330466 297538 330702 297774
rect 330146 297218 330382 297454
rect 330466 297218 330702 297454
rect 330146 263538 330382 263774
rect 330466 263538 330702 263774
rect 330146 263218 330382 263454
rect 330466 263218 330702 263454
rect 330146 229538 330382 229774
rect 330466 229538 330702 229774
rect 330146 229218 330382 229454
rect 330466 229218 330702 229454
rect 333866 711322 334102 711558
rect 334186 711322 334422 711558
rect 333866 711002 334102 711238
rect 334186 711002 334422 711238
rect 333866 675258 334102 675494
rect 334186 675258 334422 675494
rect 333866 674938 334102 675174
rect 334186 674938 334422 675174
rect 333866 641258 334102 641494
rect 334186 641258 334422 641494
rect 333866 640938 334102 641174
rect 334186 640938 334422 641174
rect 333866 607258 334102 607494
rect 334186 607258 334422 607494
rect 333866 606938 334102 607174
rect 334186 606938 334422 607174
rect 333866 573258 334102 573494
rect 334186 573258 334422 573494
rect 333866 572938 334102 573174
rect 334186 572938 334422 573174
rect 333866 539258 334102 539494
rect 334186 539258 334422 539494
rect 333866 538938 334102 539174
rect 334186 538938 334422 539174
rect 333866 505258 334102 505494
rect 334186 505258 334422 505494
rect 333866 504938 334102 505174
rect 334186 504938 334422 505174
rect 333866 471258 334102 471494
rect 334186 471258 334422 471494
rect 333866 470938 334102 471174
rect 334186 470938 334422 471174
rect 333866 437258 334102 437494
rect 334186 437258 334422 437494
rect 333866 436938 334102 437174
rect 334186 436938 334422 437174
rect 333866 403258 334102 403494
rect 334186 403258 334422 403494
rect 333866 402938 334102 403174
rect 334186 402938 334422 403174
rect 333866 369258 334102 369494
rect 334186 369258 334422 369494
rect 333866 368938 334102 369174
rect 334186 368938 334422 369174
rect 333866 335258 334102 335494
rect 334186 335258 334422 335494
rect 333866 334938 334102 335174
rect 334186 334938 334422 335174
rect 333866 301258 334102 301494
rect 334186 301258 334422 301494
rect 333866 300938 334102 301174
rect 334186 300938 334422 301174
rect 333866 267258 334102 267494
rect 334186 267258 334422 267494
rect 333866 266938 334102 267174
rect 334186 266938 334422 267174
rect 333866 233258 334102 233494
rect 334186 233258 334422 233494
rect 333866 232938 334102 233174
rect 334186 232938 334422 233174
rect 341826 704602 342062 704838
rect 342146 704602 342382 704838
rect 341826 704282 342062 704518
rect 342146 704282 342382 704518
rect 341826 683218 342062 683454
rect 342146 683218 342382 683454
rect 341826 682898 342062 683134
rect 342146 682898 342382 683134
rect 341826 649218 342062 649454
rect 342146 649218 342382 649454
rect 341826 648898 342062 649134
rect 342146 648898 342382 649134
rect 341826 615218 342062 615454
rect 342146 615218 342382 615454
rect 341826 614898 342062 615134
rect 342146 614898 342382 615134
rect 341826 581218 342062 581454
rect 342146 581218 342382 581454
rect 341826 580898 342062 581134
rect 342146 580898 342382 581134
rect 341826 547218 342062 547454
rect 342146 547218 342382 547454
rect 341826 546898 342062 547134
rect 342146 546898 342382 547134
rect 341826 513218 342062 513454
rect 342146 513218 342382 513454
rect 341826 512898 342062 513134
rect 342146 512898 342382 513134
rect 341826 479218 342062 479454
rect 342146 479218 342382 479454
rect 341826 478898 342062 479134
rect 342146 478898 342382 479134
rect 341826 445218 342062 445454
rect 342146 445218 342382 445454
rect 341826 444898 342062 445134
rect 342146 444898 342382 445134
rect 341826 411218 342062 411454
rect 342146 411218 342382 411454
rect 341826 410898 342062 411134
rect 342146 410898 342382 411134
rect 341826 377218 342062 377454
rect 342146 377218 342382 377454
rect 341826 376898 342062 377134
rect 342146 376898 342382 377134
rect 341826 343218 342062 343454
rect 342146 343218 342382 343454
rect 341826 342898 342062 343134
rect 342146 342898 342382 343134
rect 341826 309218 342062 309454
rect 342146 309218 342382 309454
rect 341826 308898 342062 309134
rect 342146 308898 342382 309134
rect 341826 275218 342062 275454
rect 342146 275218 342382 275454
rect 341826 274898 342062 275134
rect 342146 274898 342382 275134
rect 341826 241218 342062 241454
rect 342146 241218 342382 241454
rect 341826 240898 342062 241134
rect 342146 240898 342382 241134
rect 311546 210938 311782 211174
rect 311866 210938 312102 211174
rect 311546 210618 311782 210854
rect 311866 210618 312102 210854
rect 311546 176938 311782 177174
rect 311866 176938 312102 177174
rect 311546 176618 311782 176854
rect 311866 176618 312102 176854
rect 311546 142938 311782 143174
rect 311866 142938 312102 143174
rect 311546 142618 311782 142854
rect 311866 142618 312102 142854
rect 311546 108938 311782 109174
rect 311866 108938 312102 109174
rect 311546 108618 311782 108854
rect 311866 108618 312102 108854
rect 311546 74938 311782 75174
rect 311866 74938 312102 75174
rect 311546 74618 311782 74854
rect 311866 74618 312102 74854
rect 311546 40938 311782 41174
rect 311866 40938 312102 41174
rect 311546 40618 311782 40854
rect 311866 40618 312102 40854
rect 311546 6938 311782 7174
rect 311866 6938 312102 7174
rect 311546 6618 311782 6854
rect 311866 6618 312102 6854
rect 311546 -1542 311782 -1306
rect 311866 -1542 312102 -1306
rect 311546 -1862 311782 -1626
rect 311866 -1862 312102 -1626
rect 315266 180658 315502 180894
rect 315586 180658 315822 180894
rect 315266 180338 315502 180574
rect 315586 180338 315822 180574
rect 315266 146658 315502 146894
rect 315586 146658 315822 146894
rect 315266 146338 315502 146574
rect 315586 146338 315822 146574
rect 315266 112658 315502 112894
rect 315586 112658 315822 112894
rect 315266 112338 315502 112574
rect 315586 112338 315822 112574
rect 315266 78658 315502 78894
rect 315586 78658 315822 78894
rect 315266 78338 315502 78574
rect 315586 78338 315822 78574
rect 315266 44658 315502 44894
rect 315586 44658 315822 44894
rect 315266 44338 315502 44574
rect 315586 44338 315822 44574
rect 315266 10658 315502 10894
rect 315586 10658 315822 10894
rect 315266 10338 315502 10574
rect 315586 10338 315822 10574
rect 315266 -2502 315502 -2266
rect 315586 -2502 315822 -2266
rect 315266 -2822 315502 -2586
rect 315586 -2822 315822 -2586
rect 318986 184378 319222 184614
rect 319306 184378 319542 184614
rect 318986 184058 319222 184294
rect 319306 184058 319542 184294
rect 318986 150378 319222 150614
rect 319306 150378 319542 150614
rect 318986 150058 319222 150294
rect 319306 150058 319542 150294
rect 318986 116378 319222 116614
rect 319306 116378 319542 116614
rect 318986 116058 319222 116294
rect 319306 116058 319542 116294
rect 318986 82378 319222 82614
rect 319306 82378 319542 82614
rect 318986 82058 319222 82294
rect 319306 82058 319542 82294
rect 318986 48378 319222 48614
rect 319306 48378 319542 48614
rect 318986 48058 319222 48294
rect 319306 48058 319542 48294
rect 318986 14378 319222 14614
rect 319306 14378 319542 14614
rect 318986 14058 319222 14294
rect 319306 14058 319542 14294
rect 318986 -3462 319222 -3226
rect 319306 -3462 319542 -3226
rect 318986 -3782 319222 -3546
rect 319306 -3782 319542 -3546
rect 322706 188098 322942 188334
rect 323026 188098 323262 188334
rect 322706 187778 322942 188014
rect 323026 187778 323262 188014
rect 322706 154098 322942 154334
rect 323026 154098 323262 154334
rect 322706 153778 322942 154014
rect 323026 153778 323262 154014
rect 322706 120098 322942 120334
rect 323026 120098 323262 120334
rect 322706 119778 322942 120014
rect 323026 119778 323262 120014
rect 322706 86098 322942 86334
rect 323026 86098 323262 86334
rect 322706 85778 322942 86014
rect 323026 85778 323262 86014
rect 322706 52098 322942 52334
rect 323026 52098 323262 52334
rect 322706 51778 322942 52014
rect 323026 51778 323262 52014
rect 322706 18098 322942 18334
rect 323026 18098 323262 18334
rect 322706 17778 322942 18014
rect 323026 17778 323262 18014
rect 322706 -4422 322942 -4186
rect 323026 -4422 323262 -4186
rect 322706 -4742 322942 -4506
rect 323026 -4742 323262 -4506
rect 326426 191818 326662 192054
rect 326746 191818 326982 192054
rect 326426 191498 326662 191734
rect 326746 191498 326982 191734
rect 326426 157818 326662 158054
rect 326746 157818 326982 158054
rect 326426 157498 326662 157734
rect 326746 157498 326982 157734
rect 326426 123818 326662 124054
rect 326746 123818 326982 124054
rect 326426 123498 326662 123734
rect 326746 123498 326982 123734
rect 326426 89818 326662 90054
rect 326746 89818 326982 90054
rect 326426 89498 326662 89734
rect 326746 89498 326982 89734
rect 326426 55818 326662 56054
rect 326746 55818 326982 56054
rect 326426 55498 326662 55734
rect 326746 55498 326982 55734
rect 326426 21818 326662 22054
rect 326746 21818 326982 22054
rect 326426 21498 326662 21734
rect 326746 21498 326982 21734
rect 326426 -5382 326662 -5146
rect 326746 -5382 326982 -5146
rect 326426 -5702 326662 -5466
rect 326746 -5702 326982 -5466
rect 330146 195538 330382 195774
rect 330466 195538 330702 195774
rect 330146 195218 330382 195454
rect 330466 195218 330702 195454
rect 330146 161538 330382 161774
rect 330466 161538 330702 161774
rect 330146 161218 330382 161454
rect 330466 161218 330702 161454
rect 330146 127538 330382 127774
rect 330466 127538 330702 127774
rect 330146 127218 330382 127454
rect 330466 127218 330702 127454
rect 330146 93538 330382 93774
rect 330466 93538 330702 93774
rect 330146 93218 330382 93454
rect 330466 93218 330702 93454
rect 330146 59538 330382 59774
rect 330466 59538 330702 59774
rect 330146 59218 330382 59454
rect 330466 59218 330702 59454
rect 330146 25538 330382 25774
rect 330466 25538 330702 25774
rect 330146 25218 330382 25454
rect 330466 25218 330702 25454
rect 330146 -6342 330382 -6106
rect 330466 -6342 330702 -6106
rect 330146 -6662 330382 -6426
rect 330466 -6662 330702 -6426
rect 333866 199258 334102 199494
rect 334186 199258 334422 199494
rect 333866 198938 334102 199174
rect 334186 198938 334422 199174
rect 333866 165258 334102 165494
rect 334186 165258 334422 165494
rect 333866 164938 334102 165174
rect 334186 164938 334422 165174
rect 333866 131258 334102 131494
rect 334186 131258 334422 131494
rect 333866 130938 334102 131174
rect 334186 130938 334422 131174
rect 333866 97258 334102 97494
rect 334186 97258 334422 97494
rect 333866 96938 334102 97174
rect 334186 96938 334422 97174
rect 333866 63258 334102 63494
rect 334186 63258 334422 63494
rect 333866 62938 334102 63174
rect 334186 62938 334422 63174
rect 333866 29258 334102 29494
rect 334186 29258 334422 29494
rect 333866 28938 334102 29174
rect 334186 28938 334422 29174
rect 333866 -7302 334102 -7066
rect 334186 -7302 334422 -7066
rect 333866 -7622 334102 -7386
rect 334186 -7622 334422 -7386
rect 345546 705562 345782 705798
rect 345866 705562 346102 705798
rect 345546 705242 345782 705478
rect 345866 705242 346102 705478
rect 345546 686938 345782 687174
rect 345866 686938 346102 687174
rect 345546 686618 345782 686854
rect 345866 686618 346102 686854
rect 345546 652938 345782 653174
rect 345866 652938 346102 653174
rect 345546 652618 345782 652854
rect 345866 652618 346102 652854
rect 345546 618938 345782 619174
rect 345866 618938 346102 619174
rect 345546 618618 345782 618854
rect 345866 618618 346102 618854
rect 345546 584938 345782 585174
rect 345866 584938 346102 585174
rect 345546 584618 345782 584854
rect 345866 584618 346102 584854
rect 345546 550938 345782 551174
rect 345866 550938 346102 551174
rect 345546 550618 345782 550854
rect 345866 550618 346102 550854
rect 345546 516938 345782 517174
rect 345866 516938 346102 517174
rect 345546 516618 345782 516854
rect 345866 516618 346102 516854
rect 345546 482938 345782 483174
rect 345866 482938 346102 483174
rect 345546 482618 345782 482854
rect 345866 482618 346102 482854
rect 345546 448938 345782 449174
rect 345866 448938 346102 449174
rect 345546 448618 345782 448854
rect 345866 448618 346102 448854
rect 345546 414938 345782 415174
rect 345866 414938 346102 415174
rect 345546 414618 345782 414854
rect 345866 414618 346102 414854
rect 345546 380938 345782 381174
rect 345866 380938 346102 381174
rect 345546 380618 345782 380854
rect 345866 380618 346102 380854
rect 345546 346938 345782 347174
rect 345866 346938 346102 347174
rect 345546 346618 345782 346854
rect 345866 346618 346102 346854
rect 345546 312938 345782 313174
rect 345866 312938 346102 313174
rect 345546 312618 345782 312854
rect 345866 312618 346102 312854
rect 345546 278938 345782 279174
rect 345866 278938 346102 279174
rect 345546 278618 345782 278854
rect 345866 278618 346102 278854
rect 345546 244938 345782 245174
rect 345866 244938 346102 245174
rect 345546 244618 345782 244854
rect 345866 244618 346102 244854
rect 349266 706522 349502 706758
rect 349586 706522 349822 706758
rect 349266 706202 349502 706438
rect 349586 706202 349822 706438
rect 349266 690658 349502 690894
rect 349586 690658 349822 690894
rect 349266 690338 349502 690574
rect 349586 690338 349822 690574
rect 349266 656658 349502 656894
rect 349586 656658 349822 656894
rect 349266 656338 349502 656574
rect 349586 656338 349822 656574
rect 349266 622658 349502 622894
rect 349586 622658 349822 622894
rect 349266 622338 349502 622574
rect 349586 622338 349822 622574
rect 349266 588658 349502 588894
rect 349586 588658 349822 588894
rect 349266 588338 349502 588574
rect 349586 588338 349822 588574
rect 349266 554658 349502 554894
rect 349586 554658 349822 554894
rect 349266 554338 349502 554574
rect 349586 554338 349822 554574
rect 349266 520658 349502 520894
rect 349586 520658 349822 520894
rect 349266 520338 349502 520574
rect 349586 520338 349822 520574
rect 349266 486658 349502 486894
rect 349586 486658 349822 486894
rect 349266 486338 349502 486574
rect 349586 486338 349822 486574
rect 349266 452658 349502 452894
rect 349586 452658 349822 452894
rect 349266 452338 349502 452574
rect 349586 452338 349822 452574
rect 349266 418658 349502 418894
rect 349586 418658 349822 418894
rect 349266 418338 349502 418574
rect 349586 418338 349822 418574
rect 349266 384658 349502 384894
rect 349586 384658 349822 384894
rect 349266 384338 349502 384574
rect 349586 384338 349822 384574
rect 349266 350658 349502 350894
rect 349586 350658 349822 350894
rect 349266 350338 349502 350574
rect 349586 350338 349822 350574
rect 349266 316658 349502 316894
rect 349586 316658 349822 316894
rect 349266 316338 349502 316574
rect 349586 316338 349822 316574
rect 349266 282658 349502 282894
rect 349586 282658 349822 282894
rect 349266 282338 349502 282574
rect 349586 282338 349822 282574
rect 349266 248658 349502 248894
rect 349586 248658 349822 248894
rect 349266 248338 349502 248574
rect 349586 248338 349822 248574
rect 352986 707482 353222 707718
rect 353306 707482 353542 707718
rect 352986 707162 353222 707398
rect 353306 707162 353542 707398
rect 352986 694378 353222 694614
rect 353306 694378 353542 694614
rect 352986 694058 353222 694294
rect 353306 694058 353542 694294
rect 352986 660378 353222 660614
rect 353306 660378 353542 660614
rect 352986 660058 353222 660294
rect 353306 660058 353542 660294
rect 352986 626378 353222 626614
rect 353306 626378 353542 626614
rect 352986 626058 353222 626294
rect 353306 626058 353542 626294
rect 352986 592378 353222 592614
rect 353306 592378 353542 592614
rect 352986 592058 353222 592294
rect 353306 592058 353542 592294
rect 352986 558378 353222 558614
rect 353306 558378 353542 558614
rect 352986 558058 353222 558294
rect 353306 558058 353542 558294
rect 352986 524378 353222 524614
rect 353306 524378 353542 524614
rect 352986 524058 353222 524294
rect 353306 524058 353542 524294
rect 352986 490378 353222 490614
rect 353306 490378 353542 490614
rect 352986 490058 353222 490294
rect 353306 490058 353542 490294
rect 352986 456378 353222 456614
rect 353306 456378 353542 456614
rect 352986 456058 353222 456294
rect 353306 456058 353542 456294
rect 352986 422378 353222 422614
rect 353306 422378 353542 422614
rect 352986 422058 353222 422294
rect 353306 422058 353542 422294
rect 352986 388378 353222 388614
rect 353306 388378 353542 388614
rect 352986 388058 353222 388294
rect 353306 388058 353542 388294
rect 352986 354378 353222 354614
rect 353306 354378 353542 354614
rect 352986 354058 353222 354294
rect 353306 354058 353542 354294
rect 352986 320378 353222 320614
rect 353306 320378 353542 320614
rect 352986 320058 353222 320294
rect 353306 320058 353542 320294
rect 352986 286378 353222 286614
rect 353306 286378 353542 286614
rect 352986 286058 353222 286294
rect 353306 286058 353542 286294
rect 352986 252378 353222 252614
rect 353306 252378 353542 252614
rect 352986 252058 353222 252294
rect 353306 252058 353542 252294
rect 356706 708442 356942 708678
rect 357026 708442 357262 708678
rect 356706 708122 356942 708358
rect 357026 708122 357262 708358
rect 356706 698098 356942 698334
rect 357026 698098 357262 698334
rect 356706 697778 356942 698014
rect 357026 697778 357262 698014
rect 356706 664098 356942 664334
rect 357026 664098 357262 664334
rect 356706 663778 356942 664014
rect 357026 663778 357262 664014
rect 356706 630098 356942 630334
rect 357026 630098 357262 630334
rect 356706 629778 356942 630014
rect 357026 629778 357262 630014
rect 356706 596098 356942 596334
rect 357026 596098 357262 596334
rect 356706 595778 356942 596014
rect 357026 595778 357262 596014
rect 356706 562098 356942 562334
rect 357026 562098 357262 562334
rect 356706 561778 356942 562014
rect 357026 561778 357262 562014
rect 356706 528098 356942 528334
rect 357026 528098 357262 528334
rect 356706 527778 356942 528014
rect 357026 527778 357262 528014
rect 356706 494098 356942 494334
rect 357026 494098 357262 494334
rect 356706 493778 356942 494014
rect 357026 493778 357262 494014
rect 356706 460098 356942 460334
rect 357026 460098 357262 460334
rect 356706 459778 356942 460014
rect 357026 459778 357262 460014
rect 356706 426098 356942 426334
rect 357026 426098 357262 426334
rect 356706 425778 356942 426014
rect 357026 425778 357262 426014
rect 356706 392098 356942 392334
rect 357026 392098 357262 392334
rect 356706 391778 356942 392014
rect 357026 391778 357262 392014
rect 356706 358098 356942 358334
rect 357026 358098 357262 358334
rect 356706 357778 356942 358014
rect 357026 357778 357262 358014
rect 356706 324098 356942 324334
rect 357026 324098 357262 324334
rect 356706 323778 356942 324014
rect 357026 323778 357262 324014
rect 356706 290098 356942 290334
rect 357026 290098 357262 290334
rect 356706 289778 356942 290014
rect 357026 289778 357262 290014
rect 356706 256098 356942 256334
rect 357026 256098 357262 256334
rect 356706 255778 356942 256014
rect 357026 255778 357262 256014
rect 360426 709402 360662 709638
rect 360746 709402 360982 709638
rect 360426 709082 360662 709318
rect 360746 709082 360982 709318
rect 360426 667818 360662 668054
rect 360746 667818 360982 668054
rect 360426 667498 360662 667734
rect 360746 667498 360982 667734
rect 360426 633818 360662 634054
rect 360746 633818 360982 634054
rect 360426 633498 360662 633734
rect 360746 633498 360982 633734
rect 360426 599818 360662 600054
rect 360746 599818 360982 600054
rect 360426 599498 360662 599734
rect 360746 599498 360982 599734
rect 360426 565818 360662 566054
rect 360746 565818 360982 566054
rect 360426 565498 360662 565734
rect 360746 565498 360982 565734
rect 360426 531818 360662 532054
rect 360746 531818 360982 532054
rect 360426 531498 360662 531734
rect 360746 531498 360982 531734
rect 360426 497818 360662 498054
rect 360746 497818 360982 498054
rect 360426 497498 360662 497734
rect 360746 497498 360982 497734
rect 360426 463818 360662 464054
rect 360746 463818 360982 464054
rect 360426 463498 360662 463734
rect 360746 463498 360982 463734
rect 360426 429818 360662 430054
rect 360746 429818 360982 430054
rect 360426 429498 360662 429734
rect 360746 429498 360982 429734
rect 360426 395818 360662 396054
rect 360746 395818 360982 396054
rect 360426 395498 360662 395734
rect 360746 395498 360982 395734
rect 360426 361818 360662 362054
rect 360746 361818 360982 362054
rect 360426 361498 360662 361734
rect 360746 361498 360982 361734
rect 360426 327818 360662 328054
rect 360746 327818 360982 328054
rect 360426 327498 360662 327734
rect 360746 327498 360982 327734
rect 360426 293818 360662 294054
rect 360746 293818 360982 294054
rect 360426 293498 360662 293734
rect 360746 293498 360982 293734
rect 360426 259818 360662 260054
rect 360746 259818 360982 260054
rect 360426 259498 360662 259734
rect 360746 259498 360982 259734
rect 360426 225755 360662 225991
rect 360746 225755 360982 225991
rect 364146 710362 364382 710598
rect 364466 710362 364702 710598
rect 364146 710042 364382 710278
rect 364466 710042 364702 710278
rect 364146 671538 364382 671774
rect 364466 671538 364702 671774
rect 364146 671218 364382 671454
rect 364466 671218 364702 671454
rect 364146 637538 364382 637774
rect 364466 637538 364702 637774
rect 364146 637218 364382 637454
rect 364466 637218 364702 637454
rect 364146 603538 364382 603774
rect 364466 603538 364702 603774
rect 364146 603218 364382 603454
rect 364466 603218 364702 603454
rect 364146 569538 364382 569774
rect 364466 569538 364702 569774
rect 364146 569218 364382 569454
rect 364466 569218 364702 569454
rect 364146 535538 364382 535774
rect 364466 535538 364702 535774
rect 364146 535218 364382 535454
rect 364466 535218 364702 535454
rect 364146 501538 364382 501774
rect 364466 501538 364702 501774
rect 364146 501218 364382 501454
rect 364466 501218 364702 501454
rect 364146 467538 364382 467774
rect 364466 467538 364702 467774
rect 364146 467218 364382 467454
rect 364466 467218 364702 467454
rect 364146 433538 364382 433774
rect 364466 433538 364702 433774
rect 364146 433218 364382 433454
rect 364466 433218 364702 433454
rect 364146 399538 364382 399774
rect 364466 399538 364702 399774
rect 364146 399218 364382 399454
rect 364466 399218 364702 399454
rect 364146 365538 364382 365774
rect 364466 365538 364702 365774
rect 364146 365218 364382 365454
rect 364466 365218 364702 365454
rect 364146 331538 364382 331774
rect 364466 331538 364702 331774
rect 364146 331218 364382 331454
rect 364466 331218 364702 331454
rect 364146 297538 364382 297774
rect 364466 297538 364702 297774
rect 364146 297218 364382 297454
rect 364466 297218 364702 297454
rect 364146 263538 364382 263774
rect 364466 263538 364702 263774
rect 364146 263218 364382 263454
rect 364466 263218 364702 263454
rect 364146 229538 364382 229774
rect 364466 229538 364702 229774
rect 364146 229218 364382 229454
rect 364466 229218 364702 229454
rect 367866 711322 368102 711558
rect 368186 711322 368422 711558
rect 367866 711002 368102 711238
rect 368186 711002 368422 711238
rect 367866 675258 368102 675494
rect 368186 675258 368422 675494
rect 367866 674938 368102 675174
rect 368186 674938 368422 675174
rect 367866 641258 368102 641494
rect 368186 641258 368422 641494
rect 367866 640938 368102 641174
rect 368186 640938 368422 641174
rect 367866 607258 368102 607494
rect 368186 607258 368422 607494
rect 367866 606938 368102 607174
rect 368186 606938 368422 607174
rect 367866 573258 368102 573494
rect 368186 573258 368422 573494
rect 367866 572938 368102 573174
rect 368186 572938 368422 573174
rect 367866 539258 368102 539494
rect 368186 539258 368422 539494
rect 367866 538938 368102 539174
rect 368186 538938 368422 539174
rect 367866 505258 368102 505494
rect 368186 505258 368422 505494
rect 367866 504938 368102 505174
rect 368186 504938 368422 505174
rect 367866 471258 368102 471494
rect 368186 471258 368422 471494
rect 367866 470938 368102 471174
rect 368186 470938 368422 471174
rect 367866 437258 368102 437494
rect 368186 437258 368422 437494
rect 367866 436938 368102 437174
rect 368186 436938 368422 437174
rect 367866 403258 368102 403494
rect 368186 403258 368422 403494
rect 367866 402938 368102 403174
rect 368186 402938 368422 403174
rect 367866 369258 368102 369494
rect 368186 369258 368422 369494
rect 367866 368938 368102 369174
rect 368186 368938 368422 369174
rect 367866 335258 368102 335494
rect 368186 335258 368422 335494
rect 367866 334938 368102 335174
rect 368186 334938 368422 335174
rect 367866 301258 368102 301494
rect 368186 301258 368422 301494
rect 367866 300938 368102 301174
rect 368186 300938 368422 301174
rect 367866 267258 368102 267494
rect 368186 267258 368422 267494
rect 367866 266938 368102 267174
rect 368186 266938 368422 267174
rect 367866 233258 368102 233494
rect 368186 233258 368422 233494
rect 367866 232938 368102 233174
rect 368186 232938 368422 233174
rect 375826 704602 376062 704838
rect 376146 704602 376382 704838
rect 375826 704282 376062 704518
rect 376146 704282 376382 704518
rect 375826 683218 376062 683454
rect 376146 683218 376382 683454
rect 375826 682898 376062 683134
rect 376146 682898 376382 683134
rect 375826 649218 376062 649454
rect 376146 649218 376382 649454
rect 375826 648898 376062 649134
rect 376146 648898 376382 649134
rect 375826 615218 376062 615454
rect 376146 615218 376382 615454
rect 375826 614898 376062 615134
rect 376146 614898 376382 615134
rect 375826 581218 376062 581454
rect 376146 581218 376382 581454
rect 375826 580898 376062 581134
rect 376146 580898 376382 581134
rect 375826 547218 376062 547454
rect 376146 547218 376382 547454
rect 375826 546898 376062 547134
rect 376146 546898 376382 547134
rect 375826 513218 376062 513454
rect 376146 513218 376382 513454
rect 375826 512898 376062 513134
rect 376146 512898 376382 513134
rect 375826 479218 376062 479454
rect 376146 479218 376382 479454
rect 375826 478898 376062 479134
rect 376146 478898 376382 479134
rect 375826 445218 376062 445454
rect 376146 445218 376382 445454
rect 375826 444898 376062 445134
rect 376146 444898 376382 445134
rect 375826 411218 376062 411454
rect 376146 411218 376382 411454
rect 375826 410898 376062 411134
rect 376146 410898 376382 411134
rect 375826 377218 376062 377454
rect 376146 377218 376382 377454
rect 375826 376898 376062 377134
rect 376146 376898 376382 377134
rect 375826 343218 376062 343454
rect 376146 343218 376382 343454
rect 375826 342898 376062 343134
rect 376146 342898 376382 343134
rect 375826 309218 376062 309454
rect 376146 309218 376382 309454
rect 375826 308898 376062 309134
rect 376146 308898 376382 309134
rect 375826 275218 376062 275454
rect 376146 275218 376382 275454
rect 375826 274898 376062 275134
rect 376146 274898 376382 275134
rect 375826 241218 376062 241454
rect 376146 241218 376382 241454
rect 375826 240898 376062 241134
rect 376146 240898 376382 241134
rect 379546 705562 379782 705798
rect 379866 705562 380102 705798
rect 379546 705242 379782 705478
rect 379866 705242 380102 705478
rect 379546 686938 379782 687174
rect 379866 686938 380102 687174
rect 379546 686618 379782 686854
rect 379866 686618 380102 686854
rect 379546 652938 379782 653174
rect 379866 652938 380102 653174
rect 379546 652618 379782 652854
rect 379866 652618 380102 652854
rect 379546 618938 379782 619174
rect 379866 618938 380102 619174
rect 379546 618618 379782 618854
rect 379866 618618 380102 618854
rect 379546 584938 379782 585174
rect 379866 584938 380102 585174
rect 379546 584618 379782 584854
rect 379866 584618 380102 584854
rect 379546 550938 379782 551174
rect 379866 550938 380102 551174
rect 379546 550618 379782 550854
rect 379866 550618 380102 550854
rect 379546 516938 379782 517174
rect 379866 516938 380102 517174
rect 379546 516618 379782 516854
rect 379866 516618 380102 516854
rect 379546 482938 379782 483174
rect 379866 482938 380102 483174
rect 379546 482618 379782 482854
rect 379866 482618 380102 482854
rect 379546 448938 379782 449174
rect 379866 448938 380102 449174
rect 379546 448618 379782 448854
rect 379866 448618 380102 448854
rect 379546 414938 379782 415174
rect 379866 414938 380102 415174
rect 379546 414618 379782 414854
rect 379866 414618 380102 414854
rect 379546 380938 379782 381174
rect 379866 380938 380102 381174
rect 379546 380618 379782 380854
rect 379866 380618 380102 380854
rect 379546 346938 379782 347174
rect 379866 346938 380102 347174
rect 379546 346618 379782 346854
rect 379866 346618 380102 346854
rect 379546 312938 379782 313174
rect 379866 312938 380102 313174
rect 379546 312618 379782 312854
rect 379866 312618 380102 312854
rect 379546 278938 379782 279174
rect 379866 278938 380102 279174
rect 379546 278618 379782 278854
rect 379866 278618 380102 278854
rect 379546 244938 379782 245174
rect 379866 244938 380102 245174
rect 379546 244618 379782 244854
rect 379866 244618 380102 244854
rect 383266 706522 383502 706758
rect 383586 706522 383822 706758
rect 383266 706202 383502 706438
rect 383586 706202 383822 706438
rect 383266 690658 383502 690894
rect 383586 690658 383822 690894
rect 383266 690338 383502 690574
rect 383586 690338 383822 690574
rect 383266 656658 383502 656894
rect 383586 656658 383822 656894
rect 383266 656338 383502 656574
rect 383586 656338 383822 656574
rect 383266 622658 383502 622894
rect 383586 622658 383822 622894
rect 383266 622338 383502 622574
rect 383586 622338 383822 622574
rect 383266 588658 383502 588894
rect 383586 588658 383822 588894
rect 383266 588338 383502 588574
rect 383586 588338 383822 588574
rect 383266 554658 383502 554894
rect 383586 554658 383822 554894
rect 383266 554338 383502 554574
rect 383586 554338 383822 554574
rect 383266 520658 383502 520894
rect 383586 520658 383822 520894
rect 383266 520338 383502 520574
rect 383586 520338 383822 520574
rect 383266 486658 383502 486894
rect 383586 486658 383822 486894
rect 383266 486338 383502 486574
rect 383586 486338 383822 486574
rect 383266 452658 383502 452894
rect 383586 452658 383822 452894
rect 383266 452338 383502 452574
rect 383586 452338 383822 452574
rect 383266 418658 383502 418894
rect 383586 418658 383822 418894
rect 383266 418338 383502 418574
rect 383586 418338 383822 418574
rect 383266 384658 383502 384894
rect 383586 384658 383822 384894
rect 383266 384338 383502 384574
rect 383586 384338 383822 384574
rect 383266 350658 383502 350894
rect 383586 350658 383822 350894
rect 383266 350338 383502 350574
rect 383586 350338 383822 350574
rect 383266 316658 383502 316894
rect 383586 316658 383822 316894
rect 383266 316338 383502 316574
rect 383586 316338 383822 316574
rect 383266 282658 383502 282894
rect 383586 282658 383822 282894
rect 383266 282338 383502 282574
rect 383586 282338 383822 282574
rect 383266 248658 383502 248894
rect 383586 248658 383822 248894
rect 383266 248338 383502 248574
rect 383586 248338 383822 248574
rect 386986 707482 387222 707718
rect 387306 707482 387542 707718
rect 386986 707162 387222 707398
rect 387306 707162 387542 707398
rect 386986 694378 387222 694614
rect 387306 694378 387542 694614
rect 386986 694058 387222 694294
rect 387306 694058 387542 694294
rect 386986 660378 387222 660614
rect 387306 660378 387542 660614
rect 386986 660058 387222 660294
rect 387306 660058 387542 660294
rect 386986 626378 387222 626614
rect 387306 626378 387542 626614
rect 386986 626058 387222 626294
rect 387306 626058 387542 626294
rect 386986 592378 387222 592614
rect 387306 592378 387542 592614
rect 386986 592058 387222 592294
rect 387306 592058 387542 592294
rect 386986 558378 387222 558614
rect 387306 558378 387542 558614
rect 386986 558058 387222 558294
rect 387306 558058 387542 558294
rect 386986 524378 387222 524614
rect 387306 524378 387542 524614
rect 386986 524058 387222 524294
rect 387306 524058 387542 524294
rect 386986 490378 387222 490614
rect 387306 490378 387542 490614
rect 386986 490058 387222 490294
rect 387306 490058 387542 490294
rect 386986 456378 387222 456614
rect 387306 456378 387542 456614
rect 386986 456058 387222 456294
rect 387306 456058 387542 456294
rect 386986 422378 387222 422614
rect 387306 422378 387542 422614
rect 386986 422058 387222 422294
rect 387306 422058 387542 422294
rect 386986 388378 387222 388614
rect 387306 388378 387542 388614
rect 386986 388058 387222 388294
rect 387306 388058 387542 388294
rect 386986 354378 387222 354614
rect 387306 354378 387542 354614
rect 386986 354058 387222 354294
rect 387306 354058 387542 354294
rect 386986 320378 387222 320614
rect 387306 320378 387542 320614
rect 386986 320058 387222 320294
rect 387306 320058 387542 320294
rect 386986 286378 387222 286614
rect 387306 286378 387542 286614
rect 386986 286058 387222 286294
rect 387306 286058 387542 286294
rect 386986 252378 387222 252614
rect 387306 252378 387542 252614
rect 386986 252058 387222 252294
rect 387306 252058 387542 252294
rect 390706 708442 390942 708678
rect 391026 708442 391262 708678
rect 390706 708122 390942 708358
rect 391026 708122 391262 708358
rect 390706 698098 390942 698334
rect 391026 698098 391262 698334
rect 390706 697778 390942 698014
rect 391026 697778 391262 698014
rect 390706 664098 390942 664334
rect 391026 664098 391262 664334
rect 390706 663778 390942 664014
rect 391026 663778 391262 664014
rect 390706 630098 390942 630334
rect 391026 630098 391262 630334
rect 390706 629778 390942 630014
rect 391026 629778 391262 630014
rect 390706 596098 390942 596334
rect 391026 596098 391262 596334
rect 390706 595778 390942 596014
rect 391026 595778 391262 596014
rect 390706 562098 390942 562334
rect 391026 562098 391262 562334
rect 390706 561778 390942 562014
rect 391026 561778 391262 562014
rect 390706 528098 390942 528334
rect 391026 528098 391262 528334
rect 390706 527778 390942 528014
rect 391026 527778 391262 528014
rect 390706 494098 390942 494334
rect 391026 494098 391262 494334
rect 390706 493778 390942 494014
rect 391026 493778 391262 494014
rect 390706 460098 390942 460334
rect 391026 460098 391262 460334
rect 390706 459778 390942 460014
rect 391026 459778 391262 460014
rect 390706 426098 390942 426334
rect 391026 426098 391262 426334
rect 390706 425778 390942 426014
rect 391026 425778 391262 426014
rect 390706 392098 390942 392334
rect 391026 392098 391262 392334
rect 390706 391778 390942 392014
rect 391026 391778 391262 392014
rect 390706 358098 390942 358334
rect 391026 358098 391262 358334
rect 390706 357778 390942 358014
rect 391026 357778 391262 358014
rect 390706 324098 390942 324334
rect 391026 324098 391262 324334
rect 390706 323778 390942 324014
rect 391026 323778 391262 324014
rect 390706 290098 390942 290334
rect 391026 290098 391262 290334
rect 390706 289778 390942 290014
rect 391026 289778 391262 290014
rect 390706 256098 390942 256334
rect 391026 256098 391262 256334
rect 390706 255778 390942 256014
rect 391026 255778 391262 256014
rect 394426 709402 394662 709638
rect 394746 709402 394982 709638
rect 394426 709082 394662 709318
rect 394746 709082 394982 709318
rect 394426 667818 394662 668054
rect 394746 667818 394982 668054
rect 394426 667498 394662 667734
rect 394746 667498 394982 667734
rect 394426 633818 394662 634054
rect 394746 633818 394982 634054
rect 394426 633498 394662 633734
rect 394746 633498 394982 633734
rect 394426 599818 394662 600054
rect 394746 599818 394982 600054
rect 394426 599498 394662 599734
rect 394746 599498 394982 599734
rect 394426 565818 394662 566054
rect 394746 565818 394982 566054
rect 394426 565498 394662 565734
rect 394746 565498 394982 565734
rect 394426 531818 394662 532054
rect 394746 531818 394982 532054
rect 394426 531498 394662 531734
rect 394746 531498 394982 531734
rect 394426 497818 394662 498054
rect 394746 497818 394982 498054
rect 394426 497498 394662 497734
rect 394746 497498 394982 497734
rect 394426 463818 394662 464054
rect 394746 463818 394982 464054
rect 394426 463498 394662 463734
rect 394746 463498 394982 463734
rect 394426 429818 394662 430054
rect 394746 429818 394982 430054
rect 394426 429498 394662 429734
rect 394746 429498 394982 429734
rect 394426 395818 394662 396054
rect 394746 395818 394982 396054
rect 394426 395498 394662 395734
rect 394746 395498 394982 395734
rect 394426 361818 394662 362054
rect 394746 361818 394982 362054
rect 394426 361498 394662 361734
rect 394746 361498 394982 361734
rect 394426 327818 394662 328054
rect 394746 327818 394982 328054
rect 394426 327498 394662 327734
rect 394746 327498 394982 327734
rect 394426 293818 394662 294054
rect 394746 293818 394982 294054
rect 394426 293498 394662 293734
rect 394746 293498 394982 293734
rect 394426 259818 394662 260054
rect 394746 259818 394982 260054
rect 394426 259498 394662 259734
rect 394746 259498 394982 259734
rect 394426 225755 394662 225991
rect 394746 225755 394982 225991
rect 398146 710362 398382 710598
rect 398466 710362 398702 710598
rect 398146 710042 398382 710278
rect 398466 710042 398702 710278
rect 398146 671538 398382 671774
rect 398466 671538 398702 671774
rect 398146 671218 398382 671454
rect 398466 671218 398702 671454
rect 398146 637538 398382 637774
rect 398466 637538 398702 637774
rect 398146 637218 398382 637454
rect 398466 637218 398702 637454
rect 398146 603538 398382 603774
rect 398466 603538 398702 603774
rect 398146 603218 398382 603454
rect 398466 603218 398702 603454
rect 398146 569538 398382 569774
rect 398466 569538 398702 569774
rect 398146 569218 398382 569454
rect 398466 569218 398702 569454
rect 398146 535538 398382 535774
rect 398466 535538 398702 535774
rect 398146 535218 398382 535454
rect 398466 535218 398702 535454
rect 398146 501538 398382 501774
rect 398466 501538 398702 501774
rect 398146 501218 398382 501454
rect 398466 501218 398702 501454
rect 398146 467538 398382 467774
rect 398466 467538 398702 467774
rect 398146 467218 398382 467454
rect 398466 467218 398702 467454
rect 398146 433538 398382 433774
rect 398466 433538 398702 433774
rect 398146 433218 398382 433454
rect 398466 433218 398702 433454
rect 398146 399538 398382 399774
rect 398466 399538 398702 399774
rect 398146 399218 398382 399454
rect 398466 399218 398702 399454
rect 398146 365538 398382 365774
rect 398466 365538 398702 365774
rect 398146 365218 398382 365454
rect 398466 365218 398702 365454
rect 398146 331538 398382 331774
rect 398466 331538 398702 331774
rect 398146 331218 398382 331454
rect 398466 331218 398702 331454
rect 398146 297538 398382 297774
rect 398466 297538 398702 297774
rect 398146 297218 398382 297454
rect 398466 297218 398702 297454
rect 398146 263538 398382 263774
rect 398466 263538 398702 263774
rect 398146 263218 398382 263454
rect 398466 263218 398702 263454
rect 398146 229538 398382 229774
rect 398466 229538 398702 229774
rect 398146 229218 398382 229454
rect 398466 229218 398702 229454
rect 401866 711322 402102 711558
rect 402186 711322 402422 711558
rect 401866 711002 402102 711238
rect 402186 711002 402422 711238
rect 401866 675258 402102 675494
rect 402186 675258 402422 675494
rect 401866 674938 402102 675174
rect 402186 674938 402422 675174
rect 401866 641258 402102 641494
rect 402186 641258 402422 641494
rect 401866 640938 402102 641174
rect 402186 640938 402422 641174
rect 401866 607258 402102 607494
rect 402186 607258 402422 607494
rect 401866 606938 402102 607174
rect 402186 606938 402422 607174
rect 401866 573258 402102 573494
rect 402186 573258 402422 573494
rect 401866 572938 402102 573174
rect 402186 572938 402422 573174
rect 401866 539258 402102 539494
rect 402186 539258 402422 539494
rect 401866 538938 402102 539174
rect 402186 538938 402422 539174
rect 401866 505258 402102 505494
rect 402186 505258 402422 505494
rect 401866 504938 402102 505174
rect 402186 504938 402422 505174
rect 401866 471258 402102 471494
rect 402186 471258 402422 471494
rect 401866 470938 402102 471174
rect 402186 470938 402422 471174
rect 401866 437258 402102 437494
rect 402186 437258 402422 437494
rect 401866 436938 402102 437174
rect 402186 436938 402422 437174
rect 401866 403258 402102 403494
rect 402186 403258 402422 403494
rect 401866 402938 402102 403174
rect 402186 402938 402422 403174
rect 401866 369258 402102 369494
rect 402186 369258 402422 369494
rect 401866 368938 402102 369174
rect 402186 368938 402422 369174
rect 401866 335258 402102 335494
rect 402186 335258 402422 335494
rect 401866 334938 402102 335174
rect 402186 334938 402422 335174
rect 401866 301258 402102 301494
rect 402186 301258 402422 301494
rect 401866 300938 402102 301174
rect 402186 300938 402422 301174
rect 401866 267258 402102 267494
rect 402186 267258 402422 267494
rect 401866 266938 402102 267174
rect 402186 266938 402422 267174
rect 401866 233258 402102 233494
rect 402186 233258 402422 233494
rect 401866 232938 402102 233174
rect 402186 232938 402422 233174
rect 341826 207218 342062 207454
rect 342146 207218 342382 207454
rect 341826 206898 342062 207134
rect 342146 206898 342382 207134
rect 341826 173218 342062 173454
rect 342146 173218 342382 173454
rect 341826 172898 342062 173134
rect 342146 172898 342382 173134
rect 341826 139218 342062 139454
rect 342146 139218 342382 139454
rect 341826 138898 342062 139134
rect 342146 138898 342382 139134
rect 341826 105218 342062 105454
rect 342146 105218 342382 105454
rect 341826 104898 342062 105134
rect 342146 104898 342382 105134
rect 341826 71218 342062 71454
rect 342146 71218 342382 71454
rect 341826 70898 342062 71134
rect 342146 70898 342382 71134
rect 341826 37218 342062 37454
rect 342146 37218 342382 37454
rect 341826 36898 342062 37134
rect 342146 36898 342382 37134
rect 341826 3218 342062 3454
rect 342146 3218 342382 3454
rect 341826 2898 342062 3134
rect 342146 2898 342382 3134
rect 341826 -582 342062 -346
rect 342146 -582 342382 -346
rect 341826 -902 342062 -666
rect 342146 -902 342382 -666
rect 345546 210938 345782 211174
rect 345866 210938 346102 211174
rect 345546 210618 345782 210854
rect 345866 210618 346102 210854
rect 345546 176938 345782 177174
rect 345866 176938 346102 177174
rect 345546 176618 345782 176854
rect 345866 176618 346102 176854
rect 345546 142938 345782 143174
rect 345866 142938 346102 143174
rect 345546 142618 345782 142854
rect 345866 142618 346102 142854
rect 345546 108938 345782 109174
rect 345866 108938 346102 109174
rect 345546 108618 345782 108854
rect 345866 108618 346102 108854
rect 345546 74938 345782 75174
rect 345866 74938 346102 75174
rect 345546 74618 345782 74854
rect 345866 74618 346102 74854
rect 345546 40938 345782 41174
rect 345866 40938 346102 41174
rect 345546 40618 345782 40854
rect 345866 40618 346102 40854
rect 345546 6938 345782 7174
rect 345866 6938 346102 7174
rect 345546 6618 345782 6854
rect 345866 6618 346102 6854
rect 345546 -1542 345782 -1306
rect 345866 -1542 346102 -1306
rect 345546 -1862 345782 -1626
rect 345866 -1862 346102 -1626
rect 349266 180658 349502 180894
rect 349586 180658 349822 180894
rect 349266 180338 349502 180574
rect 349586 180338 349822 180574
rect 349266 146658 349502 146894
rect 349586 146658 349822 146894
rect 349266 146338 349502 146574
rect 349586 146338 349822 146574
rect 349266 112658 349502 112894
rect 349586 112658 349822 112894
rect 349266 112338 349502 112574
rect 349586 112338 349822 112574
rect 349266 78658 349502 78894
rect 349586 78658 349822 78894
rect 349266 78338 349502 78574
rect 349586 78338 349822 78574
rect 349266 44658 349502 44894
rect 349586 44658 349822 44894
rect 349266 44338 349502 44574
rect 349586 44338 349822 44574
rect 349266 10658 349502 10894
rect 349586 10658 349822 10894
rect 349266 10338 349502 10574
rect 349586 10338 349822 10574
rect 349266 -2502 349502 -2266
rect 349586 -2502 349822 -2266
rect 349266 -2822 349502 -2586
rect 349586 -2822 349822 -2586
rect 352986 184378 353222 184614
rect 353306 184378 353542 184614
rect 352986 184058 353222 184294
rect 353306 184058 353542 184294
rect 352986 150378 353222 150614
rect 353306 150378 353542 150614
rect 352986 150058 353222 150294
rect 353306 150058 353542 150294
rect 352986 116378 353222 116614
rect 353306 116378 353542 116614
rect 352986 116058 353222 116294
rect 353306 116058 353542 116294
rect 352986 82378 353222 82614
rect 353306 82378 353542 82614
rect 352986 82058 353222 82294
rect 353306 82058 353542 82294
rect 352986 48378 353222 48614
rect 353306 48378 353542 48614
rect 352986 48058 353222 48294
rect 353306 48058 353542 48294
rect 352986 14378 353222 14614
rect 353306 14378 353542 14614
rect 352986 14058 353222 14294
rect 353306 14058 353542 14294
rect 352986 -3462 353222 -3226
rect 353306 -3462 353542 -3226
rect 352986 -3782 353222 -3546
rect 353306 -3782 353542 -3546
rect 356706 188098 356942 188334
rect 357026 188098 357262 188334
rect 356706 187778 356942 188014
rect 357026 187778 357262 188014
rect 356706 154098 356942 154334
rect 357026 154098 357262 154334
rect 356706 153778 356942 154014
rect 357026 153778 357262 154014
rect 356706 120098 356942 120334
rect 357026 120098 357262 120334
rect 356706 119778 356942 120014
rect 357026 119778 357262 120014
rect 356706 86098 356942 86334
rect 357026 86098 357262 86334
rect 356706 85778 356942 86014
rect 357026 85778 357262 86014
rect 356706 52098 356942 52334
rect 357026 52098 357262 52334
rect 356706 51778 356942 52014
rect 357026 51778 357262 52014
rect 356706 18098 356942 18334
rect 357026 18098 357262 18334
rect 356706 17778 356942 18014
rect 357026 17778 357262 18014
rect 356706 -4422 356942 -4186
rect 357026 -4422 357262 -4186
rect 356706 -4742 356942 -4506
rect 357026 -4742 357262 -4506
rect 360426 191818 360662 192054
rect 360746 191818 360982 192054
rect 360426 191498 360662 191734
rect 360746 191498 360982 191734
rect 360426 157818 360662 158054
rect 360746 157818 360982 158054
rect 360426 157498 360662 157734
rect 360746 157498 360982 157734
rect 360426 123818 360662 124054
rect 360746 123818 360982 124054
rect 360426 123498 360662 123734
rect 360746 123498 360982 123734
rect 360426 89818 360662 90054
rect 360746 89818 360982 90054
rect 360426 89498 360662 89734
rect 360746 89498 360982 89734
rect 360426 55818 360662 56054
rect 360746 55818 360982 56054
rect 360426 55498 360662 55734
rect 360746 55498 360982 55734
rect 360426 21818 360662 22054
rect 360746 21818 360982 22054
rect 360426 21498 360662 21734
rect 360746 21498 360982 21734
rect 360426 -5382 360662 -5146
rect 360746 -5382 360982 -5146
rect 360426 -5702 360662 -5466
rect 360746 -5702 360982 -5466
rect 364146 195538 364382 195774
rect 364466 195538 364702 195774
rect 364146 195218 364382 195454
rect 364466 195218 364702 195454
rect 364146 161538 364382 161774
rect 364466 161538 364702 161774
rect 364146 161218 364382 161454
rect 364466 161218 364702 161454
rect 364146 127538 364382 127774
rect 364466 127538 364702 127774
rect 364146 127218 364382 127454
rect 364466 127218 364702 127454
rect 364146 93538 364382 93774
rect 364466 93538 364702 93774
rect 364146 93218 364382 93454
rect 364466 93218 364702 93454
rect 364146 59538 364382 59774
rect 364466 59538 364702 59774
rect 364146 59218 364382 59454
rect 364466 59218 364702 59454
rect 364146 25538 364382 25774
rect 364466 25538 364702 25774
rect 364146 25218 364382 25454
rect 364466 25218 364702 25454
rect 364146 -6342 364382 -6106
rect 364466 -6342 364702 -6106
rect 364146 -6662 364382 -6426
rect 364466 -6662 364702 -6426
rect 367866 199258 368102 199494
rect 368186 199258 368422 199494
rect 367866 198938 368102 199174
rect 368186 198938 368422 199174
rect 367866 165258 368102 165494
rect 368186 165258 368422 165494
rect 367866 164938 368102 165174
rect 368186 164938 368422 165174
rect 367866 131258 368102 131494
rect 368186 131258 368422 131494
rect 367866 130938 368102 131174
rect 368186 130938 368422 131174
rect 367866 97258 368102 97494
rect 368186 97258 368422 97494
rect 367866 96938 368102 97174
rect 368186 96938 368422 97174
rect 367866 63258 368102 63494
rect 368186 63258 368422 63494
rect 367866 62938 368102 63174
rect 368186 62938 368422 63174
rect 367866 29258 368102 29494
rect 368186 29258 368422 29494
rect 367866 28938 368102 29174
rect 368186 28938 368422 29174
rect 367866 -7302 368102 -7066
rect 368186 -7302 368422 -7066
rect 367866 -7622 368102 -7386
rect 368186 -7622 368422 -7386
rect 375826 207218 376062 207454
rect 376146 207218 376382 207454
rect 375826 206898 376062 207134
rect 376146 206898 376382 207134
rect 375826 173218 376062 173454
rect 376146 173218 376382 173454
rect 375826 172898 376062 173134
rect 376146 172898 376382 173134
rect 375826 139218 376062 139454
rect 376146 139218 376382 139454
rect 375826 138898 376062 139134
rect 376146 138898 376382 139134
rect 375826 105218 376062 105454
rect 376146 105218 376382 105454
rect 375826 104898 376062 105134
rect 376146 104898 376382 105134
rect 375826 71218 376062 71454
rect 376146 71218 376382 71454
rect 375826 70898 376062 71134
rect 376146 70898 376382 71134
rect 375826 37218 376062 37454
rect 376146 37218 376382 37454
rect 375826 36898 376062 37134
rect 376146 36898 376382 37134
rect 375826 3218 376062 3454
rect 376146 3218 376382 3454
rect 375826 2898 376062 3134
rect 376146 2898 376382 3134
rect 375826 -582 376062 -346
rect 376146 -582 376382 -346
rect 375826 -902 376062 -666
rect 376146 -902 376382 -666
rect 379546 210938 379782 211174
rect 379866 210938 380102 211174
rect 379546 210618 379782 210854
rect 379866 210618 380102 210854
rect 379546 176938 379782 177174
rect 379866 176938 380102 177174
rect 379546 176618 379782 176854
rect 379866 176618 380102 176854
rect 379546 142938 379782 143174
rect 379866 142938 380102 143174
rect 379546 142618 379782 142854
rect 379866 142618 380102 142854
rect 379546 108938 379782 109174
rect 379866 108938 380102 109174
rect 379546 108618 379782 108854
rect 379866 108618 380102 108854
rect 379546 74938 379782 75174
rect 379866 74938 380102 75174
rect 379546 74618 379782 74854
rect 379866 74618 380102 74854
rect 379546 40938 379782 41174
rect 379866 40938 380102 41174
rect 379546 40618 379782 40854
rect 379866 40618 380102 40854
rect 379546 6938 379782 7174
rect 379866 6938 380102 7174
rect 379546 6618 379782 6854
rect 379866 6618 380102 6854
rect 379546 -1542 379782 -1306
rect 379866 -1542 380102 -1306
rect 379546 -1862 379782 -1626
rect 379866 -1862 380102 -1626
rect 383266 180658 383502 180894
rect 383586 180658 383822 180894
rect 383266 180338 383502 180574
rect 383586 180338 383822 180574
rect 383266 146658 383502 146894
rect 383586 146658 383822 146894
rect 383266 146338 383502 146574
rect 383586 146338 383822 146574
rect 383266 112658 383502 112894
rect 383586 112658 383822 112894
rect 383266 112338 383502 112574
rect 383586 112338 383822 112574
rect 383266 78658 383502 78894
rect 383586 78658 383822 78894
rect 383266 78338 383502 78574
rect 383586 78338 383822 78574
rect 383266 44658 383502 44894
rect 383586 44658 383822 44894
rect 383266 44338 383502 44574
rect 383586 44338 383822 44574
rect 383266 10658 383502 10894
rect 383586 10658 383822 10894
rect 383266 10338 383502 10574
rect 383586 10338 383822 10574
rect 383266 -2502 383502 -2266
rect 383586 -2502 383822 -2266
rect 383266 -2822 383502 -2586
rect 383586 -2822 383822 -2586
rect 386986 184378 387222 184614
rect 387306 184378 387542 184614
rect 386986 184058 387222 184294
rect 387306 184058 387542 184294
rect 386986 150378 387222 150614
rect 387306 150378 387542 150614
rect 386986 150058 387222 150294
rect 387306 150058 387542 150294
rect 386986 116378 387222 116614
rect 387306 116378 387542 116614
rect 386986 116058 387222 116294
rect 387306 116058 387542 116294
rect 386986 82378 387222 82614
rect 387306 82378 387542 82614
rect 386986 82058 387222 82294
rect 387306 82058 387542 82294
rect 386986 48378 387222 48614
rect 387306 48378 387542 48614
rect 386986 48058 387222 48294
rect 387306 48058 387542 48294
rect 386986 14378 387222 14614
rect 387306 14378 387542 14614
rect 386986 14058 387222 14294
rect 387306 14058 387542 14294
rect 386986 -3462 387222 -3226
rect 387306 -3462 387542 -3226
rect 386986 -3782 387222 -3546
rect 387306 -3782 387542 -3546
rect 390706 188098 390942 188334
rect 391026 188098 391262 188334
rect 390706 187778 390942 188014
rect 391026 187778 391262 188014
rect 390706 154098 390942 154334
rect 391026 154098 391262 154334
rect 390706 153778 390942 154014
rect 391026 153778 391262 154014
rect 390706 120098 390942 120334
rect 391026 120098 391262 120334
rect 390706 119778 390942 120014
rect 391026 119778 391262 120014
rect 390706 86098 390942 86334
rect 391026 86098 391262 86334
rect 390706 85778 390942 86014
rect 391026 85778 391262 86014
rect 390706 52098 390942 52334
rect 391026 52098 391262 52334
rect 390706 51778 390942 52014
rect 391026 51778 391262 52014
rect 390706 18098 390942 18334
rect 391026 18098 391262 18334
rect 390706 17778 390942 18014
rect 391026 17778 391262 18014
rect 390706 -4422 390942 -4186
rect 391026 -4422 391262 -4186
rect 390706 -4742 390942 -4506
rect 391026 -4742 391262 -4506
rect 394426 191818 394662 192054
rect 394746 191818 394982 192054
rect 394426 191498 394662 191734
rect 394746 191498 394982 191734
rect 394426 157818 394662 158054
rect 394746 157818 394982 158054
rect 394426 157498 394662 157734
rect 394746 157498 394982 157734
rect 394426 123818 394662 124054
rect 394746 123818 394982 124054
rect 394426 123498 394662 123734
rect 394746 123498 394982 123734
rect 394426 89818 394662 90054
rect 394746 89818 394982 90054
rect 394426 89498 394662 89734
rect 394746 89498 394982 89734
rect 394426 55818 394662 56054
rect 394746 55818 394982 56054
rect 394426 55498 394662 55734
rect 394746 55498 394982 55734
rect 394426 21818 394662 22054
rect 394746 21818 394982 22054
rect 394426 21498 394662 21734
rect 394746 21498 394982 21734
rect 394426 -5382 394662 -5146
rect 394746 -5382 394982 -5146
rect 394426 -5702 394662 -5466
rect 394746 -5702 394982 -5466
rect 398146 195538 398382 195774
rect 398466 195538 398702 195774
rect 398146 195218 398382 195454
rect 398466 195218 398702 195454
rect 398146 161538 398382 161774
rect 398466 161538 398702 161774
rect 398146 161218 398382 161454
rect 398466 161218 398702 161454
rect 398146 127538 398382 127774
rect 398466 127538 398702 127774
rect 398146 127218 398382 127454
rect 398466 127218 398702 127454
rect 398146 93538 398382 93774
rect 398466 93538 398702 93774
rect 398146 93218 398382 93454
rect 398466 93218 398702 93454
rect 398146 59538 398382 59774
rect 398466 59538 398702 59774
rect 398146 59218 398382 59454
rect 398466 59218 398702 59454
rect 398146 25538 398382 25774
rect 398466 25538 398702 25774
rect 398146 25218 398382 25454
rect 398466 25218 398702 25454
rect 398146 -6342 398382 -6106
rect 398466 -6342 398702 -6106
rect 398146 -6662 398382 -6426
rect 398466 -6662 398702 -6426
rect 401866 199258 402102 199494
rect 402186 199258 402422 199494
rect 401866 198938 402102 199174
rect 402186 198938 402422 199174
rect 401866 165258 402102 165494
rect 402186 165258 402422 165494
rect 401866 164938 402102 165174
rect 402186 164938 402422 165174
rect 401866 131258 402102 131494
rect 402186 131258 402422 131494
rect 401866 130938 402102 131174
rect 402186 130938 402422 131174
rect 401866 97258 402102 97494
rect 402186 97258 402422 97494
rect 401866 96938 402102 97174
rect 402186 96938 402422 97174
rect 401866 63258 402102 63494
rect 402186 63258 402422 63494
rect 401866 62938 402102 63174
rect 402186 62938 402422 63174
rect 401866 29258 402102 29494
rect 402186 29258 402422 29494
rect 401866 28938 402102 29174
rect 402186 28938 402422 29174
rect 401866 -7302 402102 -7066
rect 402186 -7302 402422 -7066
rect 401866 -7622 402102 -7386
rect 402186 -7622 402422 -7386
rect 409826 704602 410062 704838
rect 410146 704602 410382 704838
rect 409826 704282 410062 704518
rect 410146 704282 410382 704518
rect 409826 683218 410062 683454
rect 410146 683218 410382 683454
rect 409826 682898 410062 683134
rect 410146 682898 410382 683134
rect 409826 649218 410062 649454
rect 410146 649218 410382 649454
rect 409826 648898 410062 649134
rect 410146 648898 410382 649134
rect 409826 615218 410062 615454
rect 410146 615218 410382 615454
rect 409826 614898 410062 615134
rect 410146 614898 410382 615134
rect 409826 581218 410062 581454
rect 410146 581218 410382 581454
rect 409826 580898 410062 581134
rect 410146 580898 410382 581134
rect 409826 547218 410062 547454
rect 410146 547218 410382 547454
rect 409826 546898 410062 547134
rect 410146 546898 410382 547134
rect 409826 513218 410062 513454
rect 410146 513218 410382 513454
rect 409826 512898 410062 513134
rect 410146 512898 410382 513134
rect 409826 479218 410062 479454
rect 410146 479218 410382 479454
rect 409826 478898 410062 479134
rect 410146 478898 410382 479134
rect 409826 445218 410062 445454
rect 410146 445218 410382 445454
rect 409826 444898 410062 445134
rect 410146 444898 410382 445134
rect 409826 411218 410062 411454
rect 410146 411218 410382 411454
rect 409826 410898 410062 411134
rect 410146 410898 410382 411134
rect 409826 377218 410062 377454
rect 410146 377218 410382 377454
rect 409826 376898 410062 377134
rect 410146 376898 410382 377134
rect 409826 343218 410062 343454
rect 410146 343218 410382 343454
rect 409826 342898 410062 343134
rect 410146 342898 410382 343134
rect 409826 309218 410062 309454
rect 410146 309218 410382 309454
rect 409826 308898 410062 309134
rect 410146 308898 410382 309134
rect 409826 275218 410062 275454
rect 410146 275218 410382 275454
rect 409826 274898 410062 275134
rect 410146 274898 410382 275134
rect 409826 241218 410062 241454
rect 410146 241218 410382 241454
rect 409826 240898 410062 241134
rect 410146 240898 410382 241134
rect 409826 207218 410062 207454
rect 410146 207218 410382 207454
rect 409826 206898 410062 207134
rect 410146 206898 410382 207134
rect 409826 173218 410062 173454
rect 410146 173218 410382 173454
rect 409826 172898 410062 173134
rect 410146 172898 410382 173134
rect 409826 139218 410062 139454
rect 410146 139218 410382 139454
rect 409826 138898 410062 139134
rect 410146 138898 410382 139134
rect 409826 105218 410062 105454
rect 410146 105218 410382 105454
rect 409826 104898 410062 105134
rect 410146 104898 410382 105134
rect 409826 71218 410062 71454
rect 410146 71218 410382 71454
rect 409826 70898 410062 71134
rect 410146 70898 410382 71134
rect 409826 37218 410062 37454
rect 410146 37218 410382 37454
rect 409826 36898 410062 37134
rect 410146 36898 410382 37134
rect 409826 3218 410062 3454
rect 410146 3218 410382 3454
rect 409826 2898 410062 3134
rect 410146 2898 410382 3134
rect 409826 -582 410062 -346
rect 410146 -582 410382 -346
rect 409826 -902 410062 -666
rect 410146 -902 410382 -666
rect 413546 705562 413782 705798
rect 413866 705562 414102 705798
rect 413546 705242 413782 705478
rect 413866 705242 414102 705478
rect 413546 686938 413782 687174
rect 413866 686938 414102 687174
rect 413546 686618 413782 686854
rect 413866 686618 414102 686854
rect 413546 652938 413782 653174
rect 413866 652938 414102 653174
rect 413546 652618 413782 652854
rect 413866 652618 414102 652854
rect 413546 618938 413782 619174
rect 413866 618938 414102 619174
rect 413546 618618 413782 618854
rect 413866 618618 414102 618854
rect 413546 584938 413782 585174
rect 413866 584938 414102 585174
rect 413546 584618 413782 584854
rect 413866 584618 414102 584854
rect 413546 550938 413782 551174
rect 413866 550938 414102 551174
rect 413546 550618 413782 550854
rect 413866 550618 414102 550854
rect 413546 516938 413782 517174
rect 413866 516938 414102 517174
rect 413546 516618 413782 516854
rect 413866 516618 414102 516854
rect 413546 482938 413782 483174
rect 413866 482938 414102 483174
rect 413546 482618 413782 482854
rect 413866 482618 414102 482854
rect 413546 448938 413782 449174
rect 413866 448938 414102 449174
rect 413546 448618 413782 448854
rect 413866 448618 414102 448854
rect 413546 414938 413782 415174
rect 413866 414938 414102 415174
rect 413546 414618 413782 414854
rect 413866 414618 414102 414854
rect 413546 380938 413782 381174
rect 413866 380938 414102 381174
rect 413546 380618 413782 380854
rect 413866 380618 414102 380854
rect 413546 346938 413782 347174
rect 413866 346938 414102 347174
rect 413546 346618 413782 346854
rect 413866 346618 414102 346854
rect 413546 312938 413782 313174
rect 413866 312938 414102 313174
rect 413546 312618 413782 312854
rect 413866 312618 414102 312854
rect 413546 278938 413782 279174
rect 413866 278938 414102 279174
rect 413546 278618 413782 278854
rect 413866 278618 414102 278854
rect 413546 244938 413782 245174
rect 413866 244938 414102 245174
rect 413546 244618 413782 244854
rect 413866 244618 414102 244854
rect 413546 210938 413782 211174
rect 413866 210938 414102 211174
rect 413546 210618 413782 210854
rect 413866 210618 414102 210854
rect 413546 176938 413782 177174
rect 413866 176938 414102 177174
rect 413546 176618 413782 176854
rect 413866 176618 414102 176854
rect 413546 142938 413782 143174
rect 413866 142938 414102 143174
rect 413546 142618 413782 142854
rect 413866 142618 414102 142854
rect 413546 108938 413782 109174
rect 413866 108938 414102 109174
rect 413546 108618 413782 108854
rect 413866 108618 414102 108854
rect 413546 74938 413782 75174
rect 413866 74938 414102 75174
rect 413546 74618 413782 74854
rect 413866 74618 414102 74854
rect 413546 40938 413782 41174
rect 413866 40938 414102 41174
rect 413546 40618 413782 40854
rect 413866 40618 414102 40854
rect 413546 6938 413782 7174
rect 413866 6938 414102 7174
rect 413546 6618 413782 6854
rect 413866 6618 414102 6854
rect 413546 -1542 413782 -1306
rect 413866 -1542 414102 -1306
rect 413546 -1862 413782 -1626
rect 413866 -1862 414102 -1626
rect 417266 706522 417502 706758
rect 417586 706522 417822 706758
rect 417266 706202 417502 706438
rect 417586 706202 417822 706438
rect 417266 690658 417502 690894
rect 417586 690658 417822 690894
rect 417266 690338 417502 690574
rect 417586 690338 417822 690574
rect 417266 656658 417502 656894
rect 417586 656658 417822 656894
rect 417266 656338 417502 656574
rect 417586 656338 417822 656574
rect 417266 622658 417502 622894
rect 417586 622658 417822 622894
rect 417266 622338 417502 622574
rect 417586 622338 417822 622574
rect 417266 588658 417502 588894
rect 417586 588658 417822 588894
rect 417266 588338 417502 588574
rect 417586 588338 417822 588574
rect 417266 554658 417502 554894
rect 417586 554658 417822 554894
rect 417266 554338 417502 554574
rect 417586 554338 417822 554574
rect 417266 520658 417502 520894
rect 417586 520658 417822 520894
rect 417266 520338 417502 520574
rect 417586 520338 417822 520574
rect 417266 486658 417502 486894
rect 417586 486658 417822 486894
rect 417266 486338 417502 486574
rect 417586 486338 417822 486574
rect 417266 452658 417502 452894
rect 417586 452658 417822 452894
rect 417266 452338 417502 452574
rect 417586 452338 417822 452574
rect 417266 418658 417502 418894
rect 417586 418658 417822 418894
rect 417266 418338 417502 418574
rect 417586 418338 417822 418574
rect 417266 384658 417502 384894
rect 417586 384658 417822 384894
rect 417266 384338 417502 384574
rect 417586 384338 417822 384574
rect 417266 350658 417502 350894
rect 417586 350658 417822 350894
rect 417266 350338 417502 350574
rect 417586 350338 417822 350574
rect 417266 316658 417502 316894
rect 417586 316658 417822 316894
rect 417266 316338 417502 316574
rect 417586 316338 417822 316574
rect 417266 282658 417502 282894
rect 417586 282658 417822 282894
rect 417266 282338 417502 282574
rect 417586 282338 417822 282574
rect 417266 248658 417502 248894
rect 417586 248658 417822 248894
rect 417266 248338 417502 248574
rect 417586 248338 417822 248574
rect 417266 214658 417502 214894
rect 417586 214658 417822 214894
rect 417266 214338 417502 214574
rect 417586 214338 417822 214574
rect 417266 180658 417502 180894
rect 417586 180658 417822 180894
rect 417266 180338 417502 180574
rect 417586 180338 417822 180574
rect 417266 146658 417502 146894
rect 417586 146658 417822 146894
rect 417266 146338 417502 146574
rect 417586 146338 417822 146574
rect 417266 112658 417502 112894
rect 417586 112658 417822 112894
rect 417266 112338 417502 112574
rect 417586 112338 417822 112574
rect 417266 78658 417502 78894
rect 417586 78658 417822 78894
rect 417266 78338 417502 78574
rect 417586 78338 417822 78574
rect 417266 44658 417502 44894
rect 417586 44658 417822 44894
rect 417266 44338 417502 44574
rect 417586 44338 417822 44574
rect 417266 10658 417502 10894
rect 417586 10658 417822 10894
rect 417266 10338 417502 10574
rect 417586 10338 417822 10574
rect 417266 -2502 417502 -2266
rect 417586 -2502 417822 -2266
rect 417266 -2822 417502 -2586
rect 417586 -2822 417822 -2586
rect 420986 707482 421222 707718
rect 421306 707482 421542 707718
rect 420986 707162 421222 707398
rect 421306 707162 421542 707398
rect 420986 694378 421222 694614
rect 421306 694378 421542 694614
rect 420986 694058 421222 694294
rect 421306 694058 421542 694294
rect 420986 660378 421222 660614
rect 421306 660378 421542 660614
rect 420986 660058 421222 660294
rect 421306 660058 421542 660294
rect 420986 626378 421222 626614
rect 421306 626378 421542 626614
rect 420986 626058 421222 626294
rect 421306 626058 421542 626294
rect 420986 592378 421222 592614
rect 421306 592378 421542 592614
rect 420986 592058 421222 592294
rect 421306 592058 421542 592294
rect 420986 558378 421222 558614
rect 421306 558378 421542 558614
rect 420986 558058 421222 558294
rect 421306 558058 421542 558294
rect 420986 524378 421222 524614
rect 421306 524378 421542 524614
rect 420986 524058 421222 524294
rect 421306 524058 421542 524294
rect 420986 490378 421222 490614
rect 421306 490378 421542 490614
rect 420986 490058 421222 490294
rect 421306 490058 421542 490294
rect 420986 456378 421222 456614
rect 421306 456378 421542 456614
rect 420986 456058 421222 456294
rect 421306 456058 421542 456294
rect 420986 422378 421222 422614
rect 421306 422378 421542 422614
rect 420986 422058 421222 422294
rect 421306 422058 421542 422294
rect 420986 388378 421222 388614
rect 421306 388378 421542 388614
rect 420986 388058 421222 388294
rect 421306 388058 421542 388294
rect 420986 354378 421222 354614
rect 421306 354378 421542 354614
rect 420986 354058 421222 354294
rect 421306 354058 421542 354294
rect 420986 320378 421222 320614
rect 421306 320378 421542 320614
rect 420986 320058 421222 320294
rect 421306 320058 421542 320294
rect 420986 286378 421222 286614
rect 421306 286378 421542 286614
rect 420986 286058 421222 286294
rect 421306 286058 421542 286294
rect 420986 252378 421222 252614
rect 421306 252378 421542 252614
rect 420986 252058 421222 252294
rect 421306 252058 421542 252294
rect 420986 218378 421222 218614
rect 421306 218378 421542 218614
rect 420986 218058 421222 218294
rect 421306 218058 421542 218294
rect 420986 184378 421222 184614
rect 421306 184378 421542 184614
rect 420986 184058 421222 184294
rect 421306 184058 421542 184294
rect 420986 150378 421222 150614
rect 421306 150378 421542 150614
rect 420986 150058 421222 150294
rect 421306 150058 421542 150294
rect 420986 116378 421222 116614
rect 421306 116378 421542 116614
rect 420986 116058 421222 116294
rect 421306 116058 421542 116294
rect 420986 82378 421222 82614
rect 421306 82378 421542 82614
rect 420986 82058 421222 82294
rect 421306 82058 421542 82294
rect 420986 48378 421222 48614
rect 421306 48378 421542 48614
rect 420986 48058 421222 48294
rect 421306 48058 421542 48294
rect 420986 14378 421222 14614
rect 421306 14378 421542 14614
rect 420986 14058 421222 14294
rect 421306 14058 421542 14294
rect 420986 -3462 421222 -3226
rect 421306 -3462 421542 -3226
rect 420986 -3782 421222 -3546
rect 421306 -3782 421542 -3546
rect 424706 708442 424942 708678
rect 425026 708442 425262 708678
rect 424706 708122 424942 708358
rect 425026 708122 425262 708358
rect 424706 698098 424942 698334
rect 425026 698098 425262 698334
rect 424706 697778 424942 698014
rect 425026 697778 425262 698014
rect 424706 664098 424942 664334
rect 425026 664098 425262 664334
rect 424706 663778 424942 664014
rect 425026 663778 425262 664014
rect 424706 630098 424942 630334
rect 425026 630098 425262 630334
rect 424706 629778 424942 630014
rect 425026 629778 425262 630014
rect 424706 596098 424942 596334
rect 425026 596098 425262 596334
rect 424706 595778 424942 596014
rect 425026 595778 425262 596014
rect 424706 562098 424942 562334
rect 425026 562098 425262 562334
rect 424706 561778 424942 562014
rect 425026 561778 425262 562014
rect 424706 528098 424942 528334
rect 425026 528098 425262 528334
rect 424706 527778 424942 528014
rect 425026 527778 425262 528014
rect 424706 494098 424942 494334
rect 425026 494098 425262 494334
rect 424706 493778 424942 494014
rect 425026 493778 425262 494014
rect 424706 460098 424942 460334
rect 425026 460098 425262 460334
rect 424706 459778 424942 460014
rect 425026 459778 425262 460014
rect 424706 426098 424942 426334
rect 425026 426098 425262 426334
rect 424706 425778 424942 426014
rect 425026 425778 425262 426014
rect 424706 392098 424942 392334
rect 425026 392098 425262 392334
rect 424706 391778 424942 392014
rect 425026 391778 425262 392014
rect 424706 358098 424942 358334
rect 425026 358098 425262 358334
rect 424706 357778 424942 358014
rect 425026 357778 425262 358014
rect 424706 324098 424942 324334
rect 425026 324098 425262 324334
rect 424706 323778 424942 324014
rect 425026 323778 425262 324014
rect 424706 290098 424942 290334
rect 425026 290098 425262 290334
rect 424706 289778 424942 290014
rect 425026 289778 425262 290014
rect 424706 256098 424942 256334
rect 425026 256098 425262 256334
rect 424706 255778 424942 256014
rect 425026 255778 425262 256014
rect 424706 222098 424942 222334
rect 425026 222098 425262 222334
rect 424706 221778 424942 222014
rect 425026 221778 425262 222014
rect 424706 188098 424942 188334
rect 425026 188098 425262 188334
rect 424706 187778 424942 188014
rect 425026 187778 425262 188014
rect 424706 154098 424942 154334
rect 425026 154098 425262 154334
rect 424706 153778 424942 154014
rect 425026 153778 425262 154014
rect 424706 120098 424942 120334
rect 425026 120098 425262 120334
rect 424706 119778 424942 120014
rect 425026 119778 425262 120014
rect 424706 86098 424942 86334
rect 425026 86098 425262 86334
rect 424706 85778 424942 86014
rect 425026 85778 425262 86014
rect 424706 52098 424942 52334
rect 425026 52098 425262 52334
rect 424706 51778 424942 52014
rect 425026 51778 425262 52014
rect 424706 18098 424942 18334
rect 425026 18098 425262 18334
rect 424706 17778 424942 18014
rect 425026 17778 425262 18014
rect 424706 -4422 424942 -4186
rect 425026 -4422 425262 -4186
rect 424706 -4742 424942 -4506
rect 425026 -4742 425262 -4506
rect 428426 709402 428662 709638
rect 428746 709402 428982 709638
rect 428426 709082 428662 709318
rect 428746 709082 428982 709318
rect 428426 667818 428662 668054
rect 428746 667818 428982 668054
rect 428426 667498 428662 667734
rect 428746 667498 428982 667734
rect 428426 633818 428662 634054
rect 428746 633818 428982 634054
rect 428426 633498 428662 633734
rect 428746 633498 428982 633734
rect 428426 599818 428662 600054
rect 428746 599818 428982 600054
rect 428426 599498 428662 599734
rect 428746 599498 428982 599734
rect 428426 565818 428662 566054
rect 428746 565818 428982 566054
rect 428426 565498 428662 565734
rect 428746 565498 428982 565734
rect 428426 531818 428662 532054
rect 428746 531818 428982 532054
rect 428426 531498 428662 531734
rect 428746 531498 428982 531734
rect 428426 497818 428662 498054
rect 428746 497818 428982 498054
rect 428426 497498 428662 497734
rect 428746 497498 428982 497734
rect 428426 463818 428662 464054
rect 428746 463818 428982 464054
rect 428426 463498 428662 463734
rect 428746 463498 428982 463734
rect 428426 429818 428662 430054
rect 428746 429818 428982 430054
rect 428426 429498 428662 429734
rect 428746 429498 428982 429734
rect 428426 395818 428662 396054
rect 428746 395818 428982 396054
rect 428426 395498 428662 395734
rect 428746 395498 428982 395734
rect 428426 361818 428662 362054
rect 428746 361818 428982 362054
rect 428426 361498 428662 361734
rect 428746 361498 428982 361734
rect 428426 327818 428662 328054
rect 428746 327818 428982 328054
rect 428426 327498 428662 327734
rect 428746 327498 428982 327734
rect 428426 293818 428662 294054
rect 428746 293818 428982 294054
rect 428426 293498 428662 293734
rect 428746 293498 428982 293734
rect 428426 259818 428662 260054
rect 428746 259818 428982 260054
rect 428426 259498 428662 259734
rect 428746 259498 428982 259734
rect 428426 225818 428662 226054
rect 428746 225818 428982 226054
rect 428426 225498 428662 225734
rect 428746 225498 428982 225734
rect 428426 191818 428662 192054
rect 428746 191818 428982 192054
rect 428426 191498 428662 191734
rect 428746 191498 428982 191734
rect 428426 157818 428662 158054
rect 428746 157818 428982 158054
rect 428426 157498 428662 157734
rect 428746 157498 428982 157734
rect 428426 123818 428662 124054
rect 428746 123818 428982 124054
rect 428426 123498 428662 123734
rect 428746 123498 428982 123734
rect 428426 89818 428662 90054
rect 428746 89818 428982 90054
rect 428426 89498 428662 89734
rect 428746 89498 428982 89734
rect 428426 55818 428662 56054
rect 428746 55818 428982 56054
rect 428426 55498 428662 55734
rect 428746 55498 428982 55734
rect 428426 21818 428662 22054
rect 428746 21818 428982 22054
rect 428426 21498 428662 21734
rect 428746 21498 428982 21734
rect 428426 -5382 428662 -5146
rect 428746 -5382 428982 -5146
rect 428426 -5702 428662 -5466
rect 428746 -5702 428982 -5466
rect 432146 710362 432382 710598
rect 432466 710362 432702 710598
rect 432146 710042 432382 710278
rect 432466 710042 432702 710278
rect 432146 671538 432382 671774
rect 432466 671538 432702 671774
rect 432146 671218 432382 671454
rect 432466 671218 432702 671454
rect 432146 637538 432382 637774
rect 432466 637538 432702 637774
rect 432146 637218 432382 637454
rect 432466 637218 432702 637454
rect 432146 603538 432382 603774
rect 432466 603538 432702 603774
rect 432146 603218 432382 603454
rect 432466 603218 432702 603454
rect 432146 569538 432382 569774
rect 432466 569538 432702 569774
rect 432146 569218 432382 569454
rect 432466 569218 432702 569454
rect 432146 535538 432382 535774
rect 432466 535538 432702 535774
rect 432146 535218 432382 535454
rect 432466 535218 432702 535454
rect 432146 501538 432382 501774
rect 432466 501538 432702 501774
rect 432146 501218 432382 501454
rect 432466 501218 432702 501454
rect 432146 467538 432382 467774
rect 432466 467538 432702 467774
rect 432146 467218 432382 467454
rect 432466 467218 432702 467454
rect 432146 433538 432382 433774
rect 432466 433538 432702 433774
rect 432146 433218 432382 433454
rect 432466 433218 432702 433454
rect 432146 399538 432382 399774
rect 432466 399538 432702 399774
rect 432146 399218 432382 399454
rect 432466 399218 432702 399454
rect 432146 365538 432382 365774
rect 432466 365538 432702 365774
rect 432146 365218 432382 365454
rect 432466 365218 432702 365454
rect 432146 331538 432382 331774
rect 432466 331538 432702 331774
rect 432146 331218 432382 331454
rect 432466 331218 432702 331454
rect 432146 297538 432382 297774
rect 432466 297538 432702 297774
rect 432146 297218 432382 297454
rect 432466 297218 432702 297454
rect 432146 263538 432382 263774
rect 432466 263538 432702 263774
rect 432146 263218 432382 263454
rect 432466 263218 432702 263454
rect 432146 229538 432382 229774
rect 432466 229538 432702 229774
rect 432146 229218 432382 229454
rect 432466 229218 432702 229454
rect 432146 195538 432382 195774
rect 432466 195538 432702 195774
rect 432146 195218 432382 195454
rect 432466 195218 432702 195454
rect 432146 161538 432382 161774
rect 432466 161538 432702 161774
rect 432146 161218 432382 161454
rect 432466 161218 432702 161454
rect 432146 127538 432382 127774
rect 432466 127538 432702 127774
rect 432146 127218 432382 127454
rect 432466 127218 432702 127454
rect 432146 93538 432382 93774
rect 432466 93538 432702 93774
rect 432146 93218 432382 93454
rect 432466 93218 432702 93454
rect 432146 59538 432382 59774
rect 432466 59538 432702 59774
rect 432146 59218 432382 59454
rect 432466 59218 432702 59454
rect 432146 25538 432382 25774
rect 432466 25538 432702 25774
rect 432146 25218 432382 25454
rect 432466 25218 432702 25454
rect 432146 -6342 432382 -6106
rect 432466 -6342 432702 -6106
rect 432146 -6662 432382 -6426
rect 432466 -6662 432702 -6426
rect 435866 711322 436102 711558
rect 436186 711322 436422 711558
rect 435866 711002 436102 711238
rect 436186 711002 436422 711238
rect 435866 675258 436102 675494
rect 436186 675258 436422 675494
rect 435866 674938 436102 675174
rect 436186 674938 436422 675174
rect 435866 641258 436102 641494
rect 436186 641258 436422 641494
rect 435866 640938 436102 641174
rect 436186 640938 436422 641174
rect 435866 607258 436102 607494
rect 436186 607258 436422 607494
rect 435866 606938 436102 607174
rect 436186 606938 436422 607174
rect 435866 573258 436102 573494
rect 436186 573258 436422 573494
rect 435866 572938 436102 573174
rect 436186 572938 436422 573174
rect 435866 539258 436102 539494
rect 436186 539258 436422 539494
rect 435866 538938 436102 539174
rect 436186 538938 436422 539174
rect 435866 505258 436102 505494
rect 436186 505258 436422 505494
rect 435866 504938 436102 505174
rect 436186 504938 436422 505174
rect 435866 471258 436102 471494
rect 436186 471258 436422 471494
rect 435866 470938 436102 471174
rect 436186 470938 436422 471174
rect 435866 437258 436102 437494
rect 436186 437258 436422 437494
rect 435866 436938 436102 437174
rect 436186 436938 436422 437174
rect 435866 403258 436102 403494
rect 436186 403258 436422 403494
rect 435866 402938 436102 403174
rect 436186 402938 436422 403174
rect 435866 369258 436102 369494
rect 436186 369258 436422 369494
rect 435866 368938 436102 369174
rect 436186 368938 436422 369174
rect 435866 335258 436102 335494
rect 436186 335258 436422 335494
rect 435866 334938 436102 335174
rect 436186 334938 436422 335174
rect 435866 301258 436102 301494
rect 436186 301258 436422 301494
rect 435866 300938 436102 301174
rect 436186 300938 436422 301174
rect 435866 267258 436102 267494
rect 436186 267258 436422 267494
rect 435866 266938 436102 267174
rect 436186 266938 436422 267174
rect 435866 233258 436102 233494
rect 436186 233258 436422 233494
rect 435866 232938 436102 233174
rect 436186 232938 436422 233174
rect 435866 199258 436102 199494
rect 436186 199258 436422 199494
rect 435866 198938 436102 199174
rect 436186 198938 436422 199174
rect 435866 165258 436102 165494
rect 436186 165258 436422 165494
rect 435866 164938 436102 165174
rect 436186 164938 436422 165174
rect 435866 131258 436102 131494
rect 436186 131258 436422 131494
rect 435866 130938 436102 131174
rect 436186 130938 436422 131174
rect 435866 97258 436102 97494
rect 436186 97258 436422 97494
rect 435866 96938 436102 97174
rect 436186 96938 436422 97174
rect 435866 63258 436102 63494
rect 436186 63258 436422 63494
rect 435866 62938 436102 63174
rect 436186 62938 436422 63174
rect 435866 29258 436102 29494
rect 436186 29258 436422 29494
rect 435866 28938 436102 29174
rect 436186 28938 436422 29174
rect 435866 -7302 436102 -7066
rect 436186 -7302 436422 -7066
rect 435866 -7622 436102 -7386
rect 436186 -7622 436422 -7386
rect 443826 704602 444062 704838
rect 444146 704602 444382 704838
rect 443826 704282 444062 704518
rect 444146 704282 444382 704518
rect 443826 683218 444062 683454
rect 444146 683218 444382 683454
rect 443826 682898 444062 683134
rect 444146 682898 444382 683134
rect 443826 649218 444062 649454
rect 444146 649218 444382 649454
rect 443826 648898 444062 649134
rect 444146 648898 444382 649134
rect 443826 615218 444062 615454
rect 444146 615218 444382 615454
rect 443826 614898 444062 615134
rect 444146 614898 444382 615134
rect 443826 581218 444062 581454
rect 444146 581218 444382 581454
rect 443826 580898 444062 581134
rect 444146 580898 444382 581134
rect 443826 547218 444062 547454
rect 444146 547218 444382 547454
rect 443826 546898 444062 547134
rect 444146 546898 444382 547134
rect 443826 513218 444062 513454
rect 444146 513218 444382 513454
rect 443826 512898 444062 513134
rect 444146 512898 444382 513134
rect 443826 479218 444062 479454
rect 444146 479218 444382 479454
rect 443826 478898 444062 479134
rect 444146 478898 444382 479134
rect 443826 445218 444062 445454
rect 444146 445218 444382 445454
rect 443826 444898 444062 445134
rect 444146 444898 444382 445134
rect 443826 411218 444062 411454
rect 444146 411218 444382 411454
rect 443826 410898 444062 411134
rect 444146 410898 444382 411134
rect 443826 377218 444062 377454
rect 444146 377218 444382 377454
rect 443826 376898 444062 377134
rect 444146 376898 444382 377134
rect 443826 343218 444062 343454
rect 444146 343218 444382 343454
rect 443826 342898 444062 343134
rect 444146 342898 444382 343134
rect 443826 309218 444062 309454
rect 444146 309218 444382 309454
rect 443826 308898 444062 309134
rect 444146 308898 444382 309134
rect 443826 275218 444062 275454
rect 444146 275218 444382 275454
rect 443826 274898 444062 275134
rect 444146 274898 444382 275134
rect 443826 241218 444062 241454
rect 444146 241218 444382 241454
rect 443826 240898 444062 241134
rect 444146 240898 444382 241134
rect 443826 207218 444062 207454
rect 444146 207218 444382 207454
rect 443826 206898 444062 207134
rect 444146 206898 444382 207134
rect 443826 173218 444062 173454
rect 444146 173218 444382 173454
rect 443826 172898 444062 173134
rect 444146 172898 444382 173134
rect 443826 139218 444062 139454
rect 444146 139218 444382 139454
rect 443826 138898 444062 139134
rect 444146 138898 444382 139134
rect 443826 105218 444062 105454
rect 444146 105218 444382 105454
rect 443826 104898 444062 105134
rect 444146 104898 444382 105134
rect 443826 71218 444062 71454
rect 444146 71218 444382 71454
rect 443826 70898 444062 71134
rect 444146 70898 444382 71134
rect 443826 37218 444062 37454
rect 444146 37218 444382 37454
rect 443826 36898 444062 37134
rect 444146 36898 444382 37134
rect 443826 3218 444062 3454
rect 444146 3218 444382 3454
rect 443826 2898 444062 3134
rect 444146 2898 444382 3134
rect 443826 -582 444062 -346
rect 444146 -582 444382 -346
rect 443826 -902 444062 -666
rect 444146 -902 444382 -666
rect 447546 705562 447782 705798
rect 447866 705562 448102 705798
rect 447546 705242 447782 705478
rect 447866 705242 448102 705478
rect 447546 686938 447782 687174
rect 447866 686938 448102 687174
rect 447546 686618 447782 686854
rect 447866 686618 448102 686854
rect 447546 652938 447782 653174
rect 447866 652938 448102 653174
rect 447546 652618 447782 652854
rect 447866 652618 448102 652854
rect 447546 618938 447782 619174
rect 447866 618938 448102 619174
rect 447546 618618 447782 618854
rect 447866 618618 448102 618854
rect 447546 584938 447782 585174
rect 447866 584938 448102 585174
rect 447546 584618 447782 584854
rect 447866 584618 448102 584854
rect 447546 550938 447782 551174
rect 447866 550938 448102 551174
rect 447546 550618 447782 550854
rect 447866 550618 448102 550854
rect 447546 516938 447782 517174
rect 447866 516938 448102 517174
rect 447546 516618 447782 516854
rect 447866 516618 448102 516854
rect 447546 482938 447782 483174
rect 447866 482938 448102 483174
rect 447546 482618 447782 482854
rect 447866 482618 448102 482854
rect 447546 448938 447782 449174
rect 447866 448938 448102 449174
rect 447546 448618 447782 448854
rect 447866 448618 448102 448854
rect 447546 414938 447782 415174
rect 447866 414938 448102 415174
rect 447546 414618 447782 414854
rect 447866 414618 448102 414854
rect 447546 380938 447782 381174
rect 447866 380938 448102 381174
rect 447546 380618 447782 380854
rect 447866 380618 448102 380854
rect 447546 346938 447782 347174
rect 447866 346938 448102 347174
rect 447546 346618 447782 346854
rect 447866 346618 448102 346854
rect 447546 312938 447782 313174
rect 447866 312938 448102 313174
rect 447546 312618 447782 312854
rect 447866 312618 448102 312854
rect 447546 278938 447782 279174
rect 447866 278938 448102 279174
rect 447546 278618 447782 278854
rect 447866 278618 448102 278854
rect 447546 244938 447782 245174
rect 447866 244938 448102 245174
rect 447546 244618 447782 244854
rect 447866 244618 448102 244854
rect 447546 210938 447782 211174
rect 447866 210938 448102 211174
rect 447546 210618 447782 210854
rect 447866 210618 448102 210854
rect 447546 176938 447782 177174
rect 447866 176938 448102 177174
rect 447546 176618 447782 176854
rect 447866 176618 448102 176854
rect 447546 142938 447782 143174
rect 447866 142938 448102 143174
rect 447546 142618 447782 142854
rect 447866 142618 448102 142854
rect 447546 108938 447782 109174
rect 447866 108938 448102 109174
rect 447546 108618 447782 108854
rect 447866 108618 448102 108854
rect 447546 74938 447782 75174
rect 447866 74938 448102 75174
rect 447546 74618 447782 74854
rect 447866 74618 448102 74854
rect 447546 40938 447782 41174
rect 447866 40938 448102 41174
rect 447546 40618 447782 40854
rect 447866 40618 448102 40854
rect 447546 6938 447782 7174
rect 447866 6938 448102 7174
rect 447546 6618 447782 6854
rect 447866 6618 448102 6854
rect 447546 -1542 447782 -1306
rect 447866 -1542 448102 -1306
rect 447546 -1862 447782 -1626
rect 447866 -1862 448102 -1626
rect 451266 706522 451502 706758
rect 451586 706522 451822 706758
rect 451266 706202 451502 706438
rect 451586 706202 451822 706438
rect 451266 690658 451502 690894
rect 451586 690658 451822 690894
rect 451266 690338 451502 690574
rect 451586 690338 451822 690574
rect 451266 656658 451502 656894
rect 451586 656658 451822 656894
rect 451266 656338 451502 656574
rect 451586 656338 451822 656574
rect 451266 622658 451502 622894
rect 451586 622658 451822 622894
rect 451266 622338 451502 622574
rect 451586 622338 451822 622574
rect 451266 588658 451502 588894
rect 451586 588658 451822 588894
rect 451266 588338 451502 588574
rect 451586 588338 451822 588574
rect 451266 554658 451502 554894
rect 451586 554658 451822 554894
rect 451266 554338 451502 554574
rect 451586 554338 451822 554574
rect 451266 520658 451502 520894
rect 451586 520658 451822 520894
rect 451266 520338 451502 520574
rect 451586 520338 451822 520574
rect 451266 486658 451502 486894
rect 451586 486658 451822 486894
rect 451266 486338 451502 486574
rect 451586 486338 451822 486574
rect 451266 452658 451502 452894
rect 451586 452658 451822 452894
rect 451266 452338 451502 452574
rect 451586 452338 451822 452574
rect 451266 418658 451502 418894
rect 451586 418658 451822 418894
rect 451266 418338 451502 418574
rect 451586 418338 451822 418574
rect 451266 384658 451502 384894
rect 451586 384658 451822 384894
rect 451266 384338 451502 384574
rect 451586 384338 451822 384574
rect 451266 350658 451502 350894
rect 451586 350658 451822 350894
rect 451266 350338 451502 350574
rect 451586 350338 451822 350574
rect 451266 316658 451502 316894
rect 451586 316658 451822 316894
rect 451266 316338 451502 316574
rect 451586 316338 451822 316574
rect 451266 282658 451502 282894
rect 451586 282658 451822 282894
rect 451266 282338 451502 282574
rect 451586 282338 451822 282574
rect 451266 248658 451502 248894
rect 451586 248658 451822 248894
rect 451266 248338 451502 248574
rect 451586 248338 451822 248574
rect 451266 214658 451502 214894
rect 451586 214658 451822 214894
rect 451266 214338 451502 214574
rect 451586 214338 451822 214574
rect 451266 180658 451502 180894
rect 451586 180658 451822 180894
rect 451266 180338 451502 180574
rect 451586 180338 451822 180574
rect 451266 146658 451502 146894
rect 451586 146658 451822 146894
rect 451266 146338 451502 146574
rect 451586 146338 451822 146574
rect 451266 112658 451502 112894
rect 451586 112658 451822 112894
rect 451266 112338 451502 112574
rect 451586 112338 451822 112574
rect 451266 78658 451502 78894
rect 451586 78658 451822 78894
rect 451266 78338 451502 78574
rect 451586 78338 451822 78574
rect 451266 44658 451502 44894
rect 451586 44658 451822 44894
rect 451266 44338 451502 44574
rect 451586 44338 451822 44574
rect 451266 10658 451502 10894
rect 451586 10658 451822 10894
rect 451266 10338 451502 10574
rect 451586 10338 451822 10574
rect 451266 -2502 451502 -2266
rect 451586 -2502 451822 -2266
rect 451266 -2822 451502 -2586
rect 451586 -2822 451822 -2586
rect 454986 707482 455222 707718
rect 455306 707482 455542 707718
rect 454986 707162 455222 707398
rect 455306 707162 455542 707398
rect 454986 694378 455222 694614
rect 455306 694378 455542 694614
rect 454986 694058 455222 694294
rect 455306 694058 455542 694294
rect 454986 660378 455222 660614
rect 455306 660378 455542 660614
rect 454986 660058 455222 660294
rect 455306 660058 455542 660294
rect 454986 626378 455222 626614
rect 455306 626378 455542 626614
rect 454986 626058 455222 626294
rect 455306 626058 455542 626294
rect 454986 592378 455222 592614
rect 455306 592378 455542 592614
rect 454986 592058 455222 592294
rect 455306 592058 455542 592294
rect 454986 558378 455222 558614
rect 455306 558378 455542 558614
rect 454986 558058 455222 558294
rect 455306 558058 455542 558294
rect 454986 524378 455222 524614
rect 455306 524378 455542 524614
rect 454986 524058 455222 524294
rect 455306 524058 455542 524294
rect 454986 490378 455222 490614
rect 455306 490378 455542 490614
rect 454986 490058 455222 490294
rect 455306 490058 455542 490294
rect 454986 456378 455222 456614
rect 455306 456378 455542 456614
rect 454986 456058 455222 456294
rect 455306 456058 455542 456294
rect 454986 422378 455222 422614
rect 455306 422378 455542 422614
rect 454986 422058 455222 422294
rect 455306 422058 455542 422294
rect 454986 388378 455222 388614
rect 455306 388378 455542 388614
rect 454986 388058 455222 388294
rect 455306 388058 455542 388294
rect 454986 354378 455222 354614
rect 455306 354378 455542 354614
rect 454986 354058 455222 354294
rect 455306 354058 455542 354294
rect 454986 320378 455222 320614
rect 455306 320378 455542 320614
rect 454986 320058 455222 320294
rect 455306 320058 455542 320294
rect 454986 286378 455222 286614
rect 455306 286378 455542 286614
rect 454986 286058 455222 286294
rect 455306 286058 455542 286294
rect 454986 252378 455222 252614
rect 455306 252378 455542 252614
rect 454986 252058 455222 252294
rect 455306 252058 455542 252294
rect 454986 218378 455222 218614
rect 455306 218378 455542 218614
rect 454986 218058 455222 218294
rect 455306 218058 455542 218294
rect 454986 184378 455222 184614
rect 455306 184378 455542 184614
rect 454986 184058 455222 184294
rect 455306 184058 455542 184294
rect 454986 150378 455222 150614
rect 455306 150378 455542 150614
rect 454986 150058 455222 150294
rect 455306 150058 455542 150294
rect 454986 116378 455222 116614
rect 455306 116378 455542 116614
rect 454986 116058 455222 116294
rect 455306 116058 455542 116294
rect 454986 82378 455222 82614
rect 455306 82378 455542 82614
rect 454986 82058 455222 82294
rect 455306 82058 455542 82294
rect 454986 48378 455222 48614
rect 455306 48378 455542 48614
rect 454986 48058 455222 48294
rect 455306 48058 455542 48294
rect 454986 14378 455222 14614
rect 455306 14378 455542 14614
rect 454986 14058 455222 14294
rect 455306 14058 455542 14294
rect 454986 -3462 455222 -3226
rect 455306 -3462 455542 -3226
rect 454986 -3782 455222 -3546
rect 455306 -3782 455542 -3546
rect 458706 708442 458942 708678
rect 459026 708442 459262 708678
rect 458706 708122 458942 708358
rect 459026 708122 459262 708358
rect 458706 698098 458942 698334
rect 459026 698098 459262 698334
rect 458706 697778 458942 698014
rect 459026 697778 459262 698014
rect 458706 664098 458942 664334
rect 459026 664098 459262 664334
rect 458706 663778 458942 664014
rect 459026 663778 459262 664014
rect 458706 630098 458942 630334
rect 459026 630098 459262 630334
rect 458706 629778 458942 630014
rect 459026 629778 459262 630014
rect 458706 596098 458942 596334
rect 459026 596098 459262 596334
rect 458706 595778 458942 596014
rect 459026 595778 459262 596014
rect 458706 562098 458942 562334
rect 459026 562098 459262 562334
rect 458706 561778 458942 562014
rect 459026 561778 459262 562014
rect 458706 528098 458942 528334
rect 459026 528098 459262 528334
rect 458706 527778 458942 528014
rect 459026 527778 459262 528014
rect 458706 494098 458942 494334
rect 459026 494098 459262 494334
rect 458706 493778 458942 494014
rect 459026 493778 459262 494014
rect 458706 460098 458942 460334
rect 459026 460098 459262 460334
rect 458706 459778 458942 460014
rect 459026 459778 459262 460014
rect 458706 426098 458942 426334
rect 459026 426098 459262 426334
rect 458706 425778 458942 426014
rect 459026 425778 459262 426014
rect 458706 392098 458942 392334
rect 459026 392098 459262 392334
rect 458706 391778 458942 392014
rect 459026 391778 459262 392014
rect 458706 358098 458942 358334
rect 459026 358098 459262 358334
rect 458706 357778 458942 358014
rect 459026 357778 459262 358014
rect 458706 324098 458942 324334
rect 459026 324098 459262 324334
rect 458706 323778 458942 324014
rect 459026 323778 459262 324014
rect 458706 290098 458942 290334
rect 459026 290098 459262 290334
rect 458706 289778 458942 290014
rect 459026 289778 459262 290014
rect 458706 256098 458942 256334
rect 459026 256098 459262 256334
rect 458706 255778 458942 256014
rect 459026 255778 459262 256014
rect 458706 222098 458942 222334
rect 459026 222098 459262 222334
rect 458706 221778 458942 222014
rect 459026 221778 459262 222014
rect 458706 188098 458942 188334
rect 459026 188098 459262 188334
rect 458706 187778 458942 188014
rect 459026 187778 459262 188014
rect 458706 154098 458942 154334
rect 459026 154098 459262 154334
rect 458706 153778 458942 154014
rect 459026 153778 459262 154014
rect 458706 120098 458942 120334
rect 459026 120098 459262 120334
rect 458706 119778 458942 120014
rect 459026 119778 459262 120014
rect 458706 86098 458942 86334
rect 459026 86098 459262 86334
rect 458706 85778 458942 86014
rect 459026 85778 459262 86014
rect 458706 52098 458942 52334
rect 459026 52098 459262 52334
rect 458706 51778 458942 52014
rect 459026 51778 459262 52014
rect 458706 18098 458942 18334
rect 459026 18098 459262 18334
rect 458706 17778 458942 18014
rect 459026 17778 459262 18014
rect 458706 -4422 458942 -4186
rect 459026 -4422 459262 -4186
rect 458706 -4742 458942 -4506
rect 459026 -4742 459262 -4506
rect 462426 709402 462662 709638
rect 462746 709402 462982 709638
rect 462426 709082 462662 709318
rect 462746 709082 462982 709318
rect 462426 667818 462662 668054
rect 462746 667818 462982 668054
rect 462426 667498 462662 667734
rect 462746 667498 462982 667734
rect 462426 633818 462662 634054
rect 462746 633818 462982 634054
rect 462426 633498 462662 633734
rect 462746 633498 462982 633734
rect 462426 599818 462662 600054
rect 462746 599818 462982 600054
rect 462426 599498 462662 599734
rect 462746 599498 462982 599734
rect 462426 565818 462662 566054
rect 462746 565818 462982 566054
rect 462426 565498 462662 565734
rect 462746 565498 462982 565734
rect 462426 531818 462662 532054
rect 462746 531818 462982 532054
rect 462426 531498 462662 531734
rect 462746 531498 462982 531734
rect 462426 497818 462662 498054
rect 462746 497818 462982 498054
rect 462426 497498 462662 497734
rect 462746 497498 462982 497734
rect 462426 463818 462662 464054
rect 462746 463818 462982 464054
rect 462426 463498 462662 463734
rect 462746 463498 462982 463734
rect 462426 429818 462662 430054
rect 462746 429818 462982 430054
rect 462426 429498 462662 429734
rect 462746 429498 462982 429734
rect 462426 395818 462662 396054
rect 462746 395818 462982 396054
rect 462426 395498 462662 395734
rect 462746 395498 462982 395734
rect 462426 361818 462662 362054
rect 462746 361818 462982 362054
rect 462426 361498 462662 361734
rect 462746 361498 462982 361734
rect 462426 327818 462662 328054
rect 462746 327818 462982 328054
rect 462426 327498 462662 327734
rect 462746 327498 462982 327734
rect 462426 293818 462662 294054
rect 462746 293818 462982 294054
rect 462426 293498 462662 293734
rect 462746 293498 462982 293734
rect 462426 259818 462662 260054
rect 462746 259818 462982 260054
rect 462426 259498 462662 259734
rect 462746 259498 462982 259734
rect 462426 225818 462662 226054
rect 462746 225818 462982 226054
rect 462426 225498 462662 225734
rect 462746 225498 462982 225734
rect 462426 191818 462662 192054
rect 462746 191818 462982 192054
rect 462426 191498 462662 191734
rect 462746 191498 462982 191734
rect 462426 157818 462662 158054
rect 462746 157818 462982 158054
rect 462426 157498 462662 157734
rect 462746 157498 462982 157734
rect 462426 123818 462662 124054
rect 462746 123818 462982 124054
rect 462426 123498 462662 123734
rect 462746 123498 462982 123734
rect 462426 89818 462662 90054
rect 462746 89818 462982 90054
rect 462426 89498 462662 89734
rect 462746 89498 462982 89734
rect 462426 55818 462662 56054
rect 462746 55818 462982 56054
rect 462426 55498 462662 55734
rect 462746 55498 462982 55734
rect 462426 21818 462662 22054
rect 462746 21818 462982 22054
rect 462426 21498 462662 21734
rect 462746 21498 462982 21734
rect 462426 -5382 462662 -5146
rect 462746 -5382 462982 -5146
rect 462426 -5702 462662 -5466
rect 462746 -5702 462982 -5466
rect 466146 710362 466382 710598
rect 466466 710362 466702 710598
rect 466146 710042 466382 710278
rect 466466 710042 466702 710278
rect 466146 671538 466382 671774
rect 466466 671538 466702 671774
rect 466146 671218 466382 671454
rect 466466 671218 466702 671454
rect 466146 637538 466382 637774
rect 466466 637538 466702 637774
rect 466146 637218 466382 637454
rect 466466 637218 466702 637454
rect 466146 603538 466382 603774
rect 466466 603538 466702 603774
rect 466146 603218 466382 603454
rect 466466 603218 466702 603454
rect 466146 569538 466382 569774
rect 466466 569538 466702 569774
rect 466146 569218 466382 569454
rect 466466 569218 466702 569454
rect 466146 535538 466382 535774
rect 466466 535538 466702 535774
rect 466146 535218 466382 535454
rect 466466 535218 466702 535454
rect 466146 501538 466382 501774
rect 466466 501538 466702 501774
rect 466146 501218 466382 501454
rect 466466 501218 466702 501454
rect 466146 467538 466382 467774
rect 466466 467538 466702 467774
rect 466146 467218 466382 467454
rect 466466 467218 466702 467454
rect 466146 433538 466382 433774
rect 466466 433538 466702 433774
rect 466146 433218 466382 433454
rect 466466 433218 466702 433454
rect 466146 399538 466382 399774
rect 466466 399538 466702 399774
rect 466146 399218 466382 399454
rect 466466 399218 466702 399454
rect 466146 365538 466382 365774
rect 466466 365538 466702 365774
rect 466146 365218 466382 365454
rect 466466 365218 466702 365454
rect 466146 331538 466382 331774
rect 466466 331538 466702 331774
rect 466146 331218 466382 331454
rect 466466 331218 466702 331454
rect 466146 297538 466382 297774
rect 466466 297538 466702 297774
rect 466146 297218 466382 297454
rect 466466 297218 466702 297454
rect 466146 263538 466382 263774
rect 466466 263538 466702 263774
rect 466146 263218 466382 263454
rect 466466 263218 466702 263454
rect 466146 229538 466382 229774
rect 466466 229538 466702 229774
rect 466146 229218 466382 229454
rect 466466 229218 466702 229454
rect 466146 195538 466382 195774
rect 466466 195538 466702 195774
rect 466146 195218 466382 195454
rect 466466 195218 466702 195454
rect 466146 161538 466382 161774
rect 466466 161538 466702 161774
rect 466146 161218 466382 161454
rect 466466 161218 466702 161454
rect 466146 127538 466382 127774
rect 466466 127538 466702 127774
rect 466146 127218 466382 127454
rect 466466 127218 466702 127454
rect 466146 93538 466382 93774
rect 466466 93538 466702 93774
rect 466146 93218 466382 93454
rect 466466 93218 466702 93454
rect 466146 59538 466382 59774
rect 466466 59538 466702 59774
rect 466146 59218 466382 59454
rect 466466 59218 466702 59454
rect 466146 25538 466382 25774
rect 466466 25538 466702 25774
rect 466146 25218 466382 25454
rect 466466 25218 466702 25454
rect 466146 -6342 466382 -6106
rect 466466 -6342 466702 -6106
rect 466146 -6662 466382 -6426
rect 466466 -6662 466702 -6426
rect 469866 711322 470102 711558
rect 470186 711322 470422 711558
rect 469866 711002 470102 711238
rect 470186 711002 470422 711238
rect 469866 675258 470102 675494
rect 470186 675258 470422 675494
rect 469866 674938 470102 675174
rect 470186 674938 470422 675174
rect 469866 641258 470102 641494
rect 470186 641258 470422 641494
rect 469866 640938 470102 641174
rect 470186 640938 470422 641174
rect 469866 607258 470102 607494
rect 470186 607258 470422 607494
rect 469866 606938 470102 607174
rect 470186 606938 470422 607174
rect 469866 573258 470102 573494
rect 470186 573258 470422 573494
rect 469866 572938 470102 573174
rect 470186 572938 470422 573174
rect 469866 539258 470102 539494
rect 470186 539258 470422 539494
rect 469866 538938 470102 539174
rect 470186 538938 470422 539174
rect 469866 505258 470102 505494
rect 470186 505258 470422 505494
rect 469866 504938 470102 505174
rect 470186 504938 470422 505174
rect 469866 471258 470102 471494
rect 470186 471258 470422 471494
rect 469866 470938 470102 471174
rect 470186 470938 470422 471174
rect 469866 437258 470102 437494
rect 470186 437258 470422 437494
rect 469866 436938 470102 437174
rect 470186 436938 470422 437174
rect 469866 403258 470102 403494
rect 470186 403258 470422 403494
rect 469866 402938 470102 403174
rect 470186 402938 470422 403174
rect 469866 369258 470102 369494
rect 470186 369258 470422 369494
rect 469866 368938 470102 369174
rect 470186 368938 470422 369174
rect 469866 335258 470102 335494
rect 470186 335258 470422 335494
rect 469866 334938 470102 335174
rect 470186 334938 470422 335174
rect 469866 301258 470102 301494
rect 470186 301258 470422 301494
rect 469866 300938 470102 301174
rect 470186 300938 470422 301174
rect 469866 267258 470102 267494
rect 470186 267258 470422 267494
rect 469866 266938 470102 267174
rect 470186 266938 470422 267174
rect 469866 233258 470102 233494
rect 470186 233258 470422 233494
rect 469866 232938 470102 233174
rect 470186 232938 470422 233174
rect 469866 199258 470102 199494
rect 470186 199258 470422 199494
rect 469866 198938 470102 199174
rect 470186 198938 470422 199174
rect 469866 165258 470102 165494
rect 470186 165258 470422 165494
rect 469866 164938 470102 165174
rect 470186 164938 470422 165174
rect 469866 131258 470102 131494
rect 470186 131258 470422 131494
rect 469866 130938 470102 131174
rect 470186 130938 470422 131174
rect 469866 97258 470102 97494
rect 470186 97258 470422 97494
rect 469866 96938 470102 97174
rect 470186 96938 470422 97174
rect 469866 63258 470102 63494
rect 470186 63258 470422 63494
rect 469866 62938 470102 63174
rect 470186 62938 470422 63174
rect 469866 29258 470102 29494
rect 470186 29258 470422 29494
rect 469866 28938 470102 29174
rect 470186 28938 470422 29174
rect 469866 -7302 470102 -7066
rect 470186 -7302 470422 -7066
rect 469866 -7622 470102 -7386
rect 470186 -7622 470422 -7386
rect 477826 704602 478062 704838
rect 478146 704602 478382 704838
rect 477826 704282 478062 704518
rect 478146 704282 478382 704518
rect 477826 683218 478062 683454
rect 478146 683218 478382 683454
rect 477826 682898 478062 683134
rect 478146 682898 478382 683134
rect 477826 649218 478062 649454
rect 478146 649218 478382 649454
rect 477826 648898 478062 649134
rect 478146 648898 478382 649134
rect 477826 615218 478062 615454
rect 478146 615218 478382 615454
rect 477826 614898 478062 615134
rect 478146 614898 478382 615134
rect 477826 581218 478062 581454
rect 478146 581218 478382 581454
rect 477826 580898 478062 581134
rect 478146 580898 478382 581134
rect 477826 547218 478062 547454
rect 478146 547218 478382 547454
rect 477826 546898 478062 547134
rect 478146 546898 478382 547134
rect 477826 513218 478062 513454
rect 478146 513218 478382 513454
rect 477826 512898 478062 513134
rect 478146 512898 478382 513134
rect 477826 479218 478062 479454
rect 478146 479218 478382 479454
rect 477826 478898 478062 479134
rect 478146 478898 478382 479134
rect 477826 445218 478062 445454
rect 478146 445218 478382 445454
rect 477826 444898 478062 445134
rect 478146 444898 478382 445134
rect 477826 411218 478062 411454
rect 478146 411218 478382 411454
rect 477826 410898 478062 411134
rect 478146 410898 478382 411134
rect 477826 377218 478062 377454
rect 478146 377218 478382 377454
rect 477826 376898 478062 377134
rect 478146 376898 478382 377134
rect 477826 343218 478062 343454
rect 478146 343218 478382 343454
rect 477826 342898 478062 343134
rect 478146 342898 478382 343134
rect 477826 309218 478062 309454
rect 478146 309218 478382 309454
rect 477826 308898 478062 309134
rect 478146 308898 478382 309134
rect 477826 275218 478062 275454
rect 478146 275218 478382 275454
rect 477826 274898 478062 275134
rect 478146 274898 478382 275134
rect 477826 241218 478062 241454
rect 478146 241218 478382 241454
rect 477826 240898 478062 241134
rect 478146 240898 478382 241134
rect 477826 207218 478062 207454
rect 478146 207218 478382 207454
rect 477826 206898 478062 207134
rect 478146 206898 478382 207134
rect 477826 173218 478062 173454
rect 478146 173218 478382 173454
rect 477826 172898 478062 173134
rect 478146 172898 478382 173134
rect 477826 139218 478062 139454
rect 478146 139218 478382 139454
rect 477826 138898 478062 139134
rect 478146 138898 478382 139134
rect 477826 105218 478062 105454
rect 478146 105218 478382 105454
rect 477826 104898 478062 105134
rect 478146 104898 478382 105134
rect 477826 71218 478062 71454
rect 478146 71218 478382 71454
rect 477826 70898 478062 71134
rect 478146 70898 478382 71134
rect 477826 37218 478062 37454
rect 478146 37218 478382 37454
rect 477826 36898 478062 37134
rect 478146 36898 478382 37134
rect 477826 3218 478062 3454
rect 478146 3218 478382 3454
rect 477826 2898 478062 3134
rect 478146 2898 478382 3134
rect 477826 -582 478062 -346
rect 478146 -582 478382 -346
rect 477826 -902 478062 -666
rect 478146 -902 478382 -666
rect 481546 705562 481782 705798
rect 481866 705562 482102 705798
rect 481546 705242 481782 705478
rect 481866 705242 482102 705478
rect 481546 686938 481782 687174
rect 481866 686938 482102 687174
rect 481546 686618 481782 686854
rect 481866 686618 482102 686854
rect 481546 652938 481782 653174
rect 481866 652938 482102 653174
rect 481546 652618 481782 652854
rect 481866 652618 482102 652854
rect 481546 618938 481782 619174
rect 481866 618938 482102 619174
rect 481546 618618 481782 618854
rect 481866 618618 482102 618854
rect 481546 584938 481782 585174
rect 481866 584938 482102 585174
rect 481546 584618 481782 584854
rect 481866 584618 482102 584854
rect 481546 550938 481782 551174
rect 481866 550938 482102 551174
rect 481546 550618 481782 550854
rect 481866 550618 482102 550854
rect 481546 516938 481782 517174
rect 481866 516938 482102 517174
rect 481546 516618 481782 516854
rect 481866 516618 482102 516854
rect 481546 482938 481782 483174
rect 481866 482938 482102 483174
rect 481546 482618 481782 482854
rect 481866 482618 482102 482854
rect 481546 448938 481782 449174
rect 481866 448938 482102 449174
rect 481546 448618 481782 448854
rect 481866 448618 482102 448854
rect 481546 414938 481782 415174
rect 481866 414938 482102 415174
rect 481546 414618 481782 414854
rect 481866 414618 482102 414854
rect 481546 380938 481782 381174
rect 481866 380938 482102 381174
rect 481546 380618 481782 380854
rect 481866 380618 482102 380854
rect 481546 346938 481782 347174
rect 481866 346938 482102 347174
rect 481546 346618 481782 346854
rect 481866 346618 482102 346854
rect 481546 312938 481782 313174
rect 481866 312938 482102 313174
rect 481546 312618 481782 312854
rect 481866 312618 482102 312854
rect 481546 278938 481782 279174
rect 481866 278938 482102 279174
rect 481546 278618 481782 278854
rect 481866 278618 482102 278854
rect 481546 244938 481782 245174
rect 481866 244938 482102 245174
rect 481546 244618 481782 244854
rect 481866 244618 482102 244854
rect 481546 210938 481782 211174
rect 481866 210938 482102 211174
rect 481546 210618 481782 210854
rect 481866 210618 482102 210854
rect 481546 176938 481782 177174
rect 481866 176938 482102 177174
rect 481546 176618 481782 176854
rect 481866 176618 482102 176854
rect 481546 142938 481782 143174
rect 481866 142938 482102 143174
rect 481546 142618 481782 142854
rect 481866 142618 482102 142854
rect 481546 108938 481782 109174
rect 481866 108938 482102 109174
rect 481546 108618 481782 108854
rect 481866 108618 482102 108854
rect 481546 74938 481782 75174
rect 481866 74938 482102 75174
rect 481546 74618 481782 74854
rect 481866 74618 482102 74854
rect 481546 40938 481782 41174
rect 481866 40938 482102 41174
rect 481546 40618 481782 40854
rect 481866 40618 482102 40854
rect 481546 6938 481782 7174
rect 481866 6938 482102 7174
rect 481546 6618 481782 6854
rect 481866 6618 482102 6854
rect 481546 -1542 481782 -1306
rect 481866 -1542 482102 -1306
rect 481546 -1862 481782 -1626
rect 481866 -1862 482102 -1626
rect 485266 706522 485502 706758
rect 485586 706522 485822 706758
rect 485266 706202 485502 706438
rect 485586 706202 485822 706438
rect 485266 690658 485502 690894
rect 485586 690658 485822 690894
rect 485266 690338 485502 690574
rect 485586 690338 485822 690574
rect 485266 656658 485502 656894
rect 485586 656658 485822 656894
rect 485266 656338 485502 656574
rect 485586 656338 485822 656574
rect 485266 622658 485502 622894
rect 485586 622658 485822 622894
rect 485266 622338 485502 622574
rect 485586 622338 485822 622574
rect 485266 588658 485502 588894
rect 485586 588658 485822 588894
rect 485266 588338 485502 588574
rect 485586 588338 485822 588574
rect 485266 554658 485502 554894
rect 485586 554658 485822 554894
rect 485266 554338 485502 554574
rect 485586 554338 485822 554574
rect 485266 520658 485502 520894
rect 485586 520658 485822 520894
rect 485266 520338 485502 520574
rect 485586 520338 485822 520574
rect 485266 486658 485502 486894
rect 485586 486658 485822 486894
rect 485266 486338 485502 486574
rect 485586 486338 485822 486574
rect 485266 452658 485502 452894
rect 485586 452658 485822 452894
rect 485266 452338 485502 452574
rect 485586 452338 485822 452574
rect 485266 418658 485502 418894
rect 485586 418658 485822 418894
rect 485266 418338 485502 418574
rect 485586 418338 485822 418574
rect 485266 384658 485502 384894
rect 485586 384658 485822 384894
rect 485266 384338 485502 384574
rect 485586 384338 485822 384574
rect 485266 350658 485502 350894
rect 485586 350658 485822 350894
rect 485266 350338 485502 350574
rect 485586 350338 485822 350574
rect 485266 316658 485502 316894
rect 485586 316658 485822 316894
rect 485266 316338 485502 316574
rect 485586 316338 485822 316574
rect 485266 282658 485502 282894
rect 485586 282658 485822 282894
rect 485266 282338 485502 282574
rect 485586 282338 485822 282574
rect 485266 248658 485502 248894
rect 485586 248658 485822 248894
rect 485266 248338 485502 248574
rect 485586 248338 485822 248574
rect 485266 214658 485502 214894
rect 485586 214658 485822 214894
rect 485266 214338 485502 214574
rect 485586 214338 485822 214574
rect 485266 180658 485502 180894
rect 485586 180658 485822 180894
rect 485266 180338 485502 180574
rect 485586 180338 485822 180574
rect 485266 146658 485502 146894
rect 485586 146658 485822 146894
rect 485266 146338 485502 146574
rect 485586 146338 485822 146574
rect 485266 112658 485502 112894
rect 485586 112658 485822 112894
rect 485266 112338 485502 112574
rect 485586 112338 485822 112574
rect 485266 78658 485502 78894
rect 485586 78658 485822 78894
rect 485266 78338 485502 78574
rect 485586 78338 485822 78574
rect 485266 44658 485502 44894
rect 485586 44658 485822 44894
rect 485266 44338 485502 44574
rect 485586 44338 485822 44574
rect 485266 10658 485502 10894
rect 485586 10658 485822 10894
rect 485266 10338 485502 10574
rect 485586 10338 485822 10574
rect 485266 -2502 485502 -2266
rect 485586 -2502 485822 -2266
rect 485266 -2822 485502 -2586
rect 485586 -2822 485822 -2586
rect 488986 707482 489222 707718
rect 489306 707482 489542 707718
rect 488986 707162 489222 707398
rect 489306 707162 489542 707398
rect 488986 694378 489222 694614
rect 489306 694378 489542 694614
rect 488986 694058 489222 694294
rect 489306 694058 489542 694294
rect 488986 660378 489222 660614
rect 489306 660378 489542 660614
rect 488986 660058 489222 660294
rect 489306 660058 489542 660294
rect 488986 626378 489222 626614
rect 489306 626378 489542 626614
rect 488986 626058 489222 626294
rect 489306 626058 489542 626294
rect 488986 592378 489222 592614
rect 489306 592378 489542 592614
rect 488986 592058 489222 592294
rect 489306 592058 489542 592294
rect 488986 558378 489222 558614
rect 489306 558378 489542 558614
rect 488986 558058 489222 558294
rect 489306 558058 489542 558294
rect 488986 524378 489222 524614
rect 489306 524378 489542 524614
rect 488986 524058 489222 524294
rect 489306 524058 489542 524294
rect 488986 490378 489222 490614
rect 489306 490378 489542 490614
rect 488986 490058 489222 490294
rect 489306 490058 489542 490294
rect 488986 456378 489222 456614
rect 489306 456378 489542 456614
rect 488986 456058 489222 456294
rect 489306 456058 489542 456294
rect 488986 422378 489222 422614
rect 489306 422378 489542 422614
rect 488986 422058 489222 422294
rect 489306 422058 489542 422294
rect 488986 388378 489222 388614
rect 489306 388378 489542 388614
rect 488986 388058 489222 388294
rect 489306 388058 489542 388294
rect 488986 354378 489222 354614
rect 489306 354378 489542 354614
rect 488986 354058 489222 354294
rect 489306 354058 489542 354294
rect 488986 320378 489222 320614
rect 489306 320378 489542 320614
rect 488986 320058 489222 320294
rect 489306 320058 489542 320294
rect 488986 286378 489222 286614
rect 489306 286378 489542 286614
rect 488986 286058 489222 286294
rect 489306 286058 489542 286294
rect 488986 252378 489222 252614
rect 489306 252378 489542 252614
rect 488986 252058 489222 252294
rect 489306 252058 489542 252294
rect 488986 218378 489222 218614
rect 489306 218378 489542 218614
rect 488986 218058 489222 218294
rect 489306 218058 489542 218294
rect 488986 184378 489222 184614
rect 489306 184378 489542 184614
rect 488986 184058 489222 184294
rect 489306 184058 489542 184294
rect 488986 150378 489222 150614
rect 489306 150378 489542 150614
rect 488986 150058 489222 150294
rect 489306 150058 489542 150294
rect 488986 116378 489222 116614
rect 489306 116378 489542 116614
rect 488986 116058 489222 116294
rect 489306 116058 489542 116294
rect 488986 82378 489222 82614
rect 489306 82378 489542 82614
rect 488986 82058 489222 82294
rect 489306 82058 489542 82294
rect 488986 48378 489222 48614
rect 489306 48378 489542 48614
rect 488986 48058 489222 48294
rect 489306 48058 489542 48294
rect 488986 14378 489222 14614
rect 489306 14378 489542 14614
rect 488986 14058 489222 14294
rect 489306 14058 489542 14294
rect 488986 -3462 489222 -3226
rect 489306 -3462 489542 -3226
rect 488986 -3782 489222 -3546
rect 489306 -3782 489542 -3546
rect 492706 708442 492942 708678
rect 493026 708442 493262 708678
rect 492706 708122 492942 708358
rect 493026 708122 493262 708358
rect 492706 698098 492942 698334
rect 493026 698098 493262 698334
rect 492706 697778 492942 698014
rect 493026 697778 493262 698014
rect 492706 664098 492942 664334
rect 493026 664098 493262 664334
rect 492706 663778 492942 664014
rect 493026 663778 493262 664014
rect 492706 630098 492942 630334
rect 493026 630098 493262 630334
rect 492706 629778 492942 630014
rect 493026 629778 493262 630014
rect 492706 596098 492942 596334
rect 493026 596098 493262 596334
rect 492706 595778 492942 596014
rect 493026 595778 493262 596014
rect 492706 562098 492942 562334
rect 493026 562098 493262 562334
rect 492706 561778 492942 562014
rect 493026 561778 493262 562014
rect 492706 528098 492942 528334
rect 493026 528098 493262 528334
rect 492706 527778 492942 528014
rect 493026 527778 493262 528014
rect 492706 494098 492942 494334
rect 493026 494098 493262 494334
rect 492706 493778 492942 494014
rect 493026 493778 493262 494014
rect 492706 460098 492942 460334
rect 493026 460098 493262 460334
rect 492706 459778 492942 460014
rect 493026 459778 493262 460014
rect 492706 426098 492942 426334
rect 493026 426098 493262 426334
rect 492706 425778 492942 426014
rect 493026 425778 493262 426014
rect 492706 392098 492942 392334
rect 493026 392098 493262 392334
rect 492706 391778 492942 392014
rect 493026 391778 493262 392014
rect 492706 358098 492942 358334
rect 493026 358098 493262 358334
rect 492706 357778 492942 358014
rect 493026 357778 493262 358014
rect 492706 324098 492942 324334
rect 493026 324098 493262 324334
rect 492706 323778 492942 324014
rect 493026 323778 493262 324014
rect 492706 290098 492942 290334
rect 493026 290098 493262 290334
rect 492706 289778 492942 290014
rect 493026 289778 493262 290014
rect 492706 256098 492942 256334
rect 493026 256098 493262 256334
rect 492706 255778 492942 256014
rect 493026 255778 493262 256014
rect 492706 222098 492942 222334
rect 493026 222098 493262 222334
rect 492706 221778 492942 222014
rect 493026 221778 493262 222014
rect 492706 188098 492942 188334
rect 493026 188098 493262 188334
rect 492706 187778 492942 188014
rect 493026 187778 493262 188014
rect 492706 154098 492942 154334
rect 493026 154098 493262 154334
rect 492706 153778 492942 154014
rect 493026 153778 493262 154014
rect 492706 120098 492942 120334
rect 493026 120098 493262 120334
rect 492706 119778 492942 120014
rect 493026 119778 493262 120014
rect 492706 86098 492942 86334
rect 493026 86098 493262 86334
rect 492706 85778 492942 86014
rect 493026 85778 493262 86014
rect 492706 52098 492942 52334
rect 493026 52098 493262 52334
rect 492706 51778 492942 52014
rect 493026 51778 493262 52014
rect 492706 18098 492942 18334
rect 493026 18098 493262 18334
rect 492706 17778 492942 18014
rect 493026 17778 493262 18014
rect 492706 -4422 492942 -4186
rect 493026 -4422 493262 -4186
rect 492706 -4742 492942 -4506
rect 493026 -4742 493262 -4506
rect 496426 709402 496662 709638
rect 496746 709402 496982 709638
rect 496426 709082 496662 709318
rect 496746 709082 496982 709318
rect 496426 667818 496662 668054
rect 496746 667818 496982 668054
rect 496426 667498 496662 667734
rect 496746 667498 496982 667734
rect 496426 633818 496662 634054
rect 496746 633818 496982 634054
rect 496426 633498 496662 633734
rect 496746 633498 496982 633734
rect 496426 599818 496662 600054
rect 496746 599818 496982 600054
rect 496426 599498 496662 599734
rect 496746 599498 496982 599734
rect 496426 565818 496662 566054
rect 496746 565818 496982 566054
rect 496426 565498 496662 565734
rect 496746 565498 496982 565734
rect 496426 531818 496662 532054
rect 496746 531818 496982 532054
rect 496426 531498 496662 531734
rect 496746 531498 496982 531734
rect 496426 497818 496662 498054
rect 496746 497818 496982 498054
rect 496426 497498 496662 497734
rect 496746 497498 496982 497734
rect 496426 463818 496662 464054
rect 496746 463818 496982 464054
rect 496426 463498 496662 463734
rect 496746 463498 496982 463734
rect 496426 429818 496662 430054
rect 496746 429818 496982 430054
rect 496426 429498 496662 429734
rect 496746 429498 496982 429734
rect 496426 395818 496662 396054
rect 496746 395818 496982 396054
rect 496426 395498 496662 395734
rect 496746 395498 496982 395734
rect 496426 361818 496662 362054
rect 496746 361818 496982 362054
rect 496426 361498 496662 361734
rect 496746 361498 496982 361734
rect 496426 327818 496662 328054
rect 496746 327818 496982 328054
rect 496426 327498 496662 327734
rect 496746 327498 496982 327734
rect 496426 293818 496662 294054
rect 496746 293818 496982 294054
rect 496426 293498 496662 293734
rect 496746 293498 496982 293734
rect 496426 259818 496662 260054
rect 496746 259818 496982 260054
rect 496426 259498 496662 259734
rect 496746 259498 496982 259734
rect 496426 225818 496662 226054
rect 496746 225818 496982 226054
rect 496426 225498 496662 225734
rect 496746 225498 496982 225734
rect 496426 191818 496662 192054
rect 496746 191818 496982 192054
rect 496426 191498 496662 191734
rect 496746 191498 496982 191734
rect 496426 157818 496662 158054
rect 496746 157818 496982 158054
rect 496426 157498 496662 157734
rect 496746 157498 496982 157734
rect 496426 123818 496662 124054
rect 496746 123818 496982 124054
rect 496426 123498 496662 123734
rect 496746 123498 496982 123734
rect 496426 89818 496662 90054
rect 496746 89818 496982 90054
rect 496426 89498 496662 89734
rect 496746 89498 496982 89734
rect 496426 55818 496662 56054
rect 496746 55818 496982 56054
rect 496426 55498 496662 55734
rect 496746 55498 496982 55734
rect 496426 21818 496662 22054
rect 496746 21818 496982 22054
rect 496426 21498 496662 21734
rect 496746 21498 496982 21734
rect 496426 -5382 496662 -5146
rect 496746 -5382 496982 -5146
rect 496426 -5702 496662 -5466
rect 496746 -5702 496982 -5466
rect 500146 710362 500382 710598
rect 500466 710362 500702 710598
rect 500146 710042 500382 710278
rect 500466 710042 500702 710278
rect 500146 671538 500382 671774
rect 500466 671538 500702 671774
rect 500146 671218 500382 671454
rect 500466 671218 500702 671454
rect 500146 637538 500382 637774
rect 500466 637538 500702 637774
rect 500146 637218 500382 637454
rect 500466 637218 500702 637454
rect 500146 603538 500382 603774
rect 500466 603538 500702 603774
rect 500146 603218 500382 603454
rect 500466 603218 500702 603454
rect 500146 569538 500382 569774
rect 500466 569538 500702 569774
rect 500146 569218 500382 569454
rect 500466 569218 500702 569454
rect 500146 535538 500382 535774
rect 500466 535538 500702 535774
rect 500146 535218 500382 535454
rect 500466 535218 500702 535454
rect 500146 501538 500382 501774
rect 500466 501538 500702 501774
rect 500146 501218 500382 501454
rect 500466 501218 500702 501454
rect 500146 467538 500382 467774
rect 500466 467538 500702 467774
rect 500146 467218 500382 467454
rect 500466 467218 500702 467454
rect 500146 433538 500382 433774
rect 500466 433538 500702 433774
rect 500146 433218 500382 433454
rect 500466 433218 500702 433454
rect 500146 399538 500382 399774
rect 500466 399538 500702 399774
rect 500146 399218 500382 399454
rect 500466 399218 500702 399454
rect 500146 365538 500382 365774
rect 500466 365538 500702 365774
rect 500146 365218 500382 365454
rect 500466 365218 500702 365454
rect 500146 331538 500382 331774
rect 500466 331538 500702 331774
rect 500146 331218 500382 331454
rect 500466 331218 500702 331454
rect 500146 297538 500382 297774
rect 500466 297538 500702 297774
rect 500146 297218 500382 297454
rect 500466 297218 500702 297454
rect 500146 263538 500382 263774
rect 500466 263538 500702 263774
rect 500146 263218 500382 263454
rect 500466 263218 500702 263454
rect 500146 229538 500382 229774
rect 500466 229538 500702 229774
rect 500146 229218 500382 229454
rect 500466 229218 500702 229454
rect 500146 195538 500382 195774
rect 500466 195538 500702 195774
rect 500146 195218 500382 195454
rect 500466 195218 500702 195454
rect 500146 161538 500382 161774
rect 500466 161538 500702 161774
rect 500146 161218 500382 161454
rect 500466 161218 500702 161454
rect 500146 127538 500382 127774
rect 500466 127538 500702 127774
rect 500146 127218 500382 127454
rect 500466 127218 500702 127454
rect 500146 93538 500382 93774
rect 500466 93538 500702 93774
rect 500146 93218 500382 93454
rect 500466 93218 500702 93454
rect 500146 59538 500382 59774
rect 500466 59538 500702 59774
rect 500146 59218 500382 59454
rect 500466 59218 500702 59454
rect 500146 25538 500382 25774
rect 500466 25538 500702 25774
rect 500146 25218 500382 25454
rect 500466 25218 500702 25454
rect 500146 -6342 500382 -6106
rect 500466 -6342 500702 -6106
rect 500146 -6662 500382 -6426
rect 500466 -6662 500702 -6426
rect 503866 711322 504102 711558
rect 504186 711322 504422 711558
rect 503866 711002 504102 711238
rect 504186 711002 504422 711238
rect 503866 675258 504102 675494
rect 504186 675258 504422 675494
rect 503866 674938 504102 675174
rect 504186 674938 504422 675174
rect 503866 641258 504102 641494
rect 504186 641258 504422 641494
rect 503866 640938 504102 641174
rect 504186 640938 504422 641174
rect 503866 607258 504102 607494
rect 504186 607258 504422 607494
rect 503866 606938 504102 607174
rect 504186 606938 504422 607174
rect 503866 573258 504102 573494
rect 504186 573258 504422 573494
rect 503866 572938 504102 573174
rect 504186 572938 504422 573174
rect 503866 539258 504102 539494
rect 504186 539258 504422 539494
rect 503866 538938 504102 539174
rect 504186 538938 504422 539174
rect 503866 505258 504102 505494
rect 504186 505258 504422 505494
rect 503866 504938 504102 505174
rect 504186 504938 504422 505174
rect 503866 471258 504102 471494
rect 504186 471258 504422 471494
rect 503866 470938 504102 471174
rect 504186 470938 504422 471174
rect 503866 437258 504102 437494
rect 504186 437258 504422 437494
rect 503866 436938 504102 437174
rect 504186 436938 504422 437174
rect 503866 403258 504102 403494
rect 504186 403258 504422 403494
rect 503866 402938 504102 403174
rect 504186 402938 504422 403174
rect 503866 369258 504102 369494
rect 504186 369258 504422 369494
rect 503866 368938 504102 369174
rect 504186 368938 504422 369174
rect 503866 335258 504102 335494
rect 504186 335258 504422 335494
rect 503866 334938 504102 335174
rect 504186 334938 504422 335174
rect 503866 301258 504102 301494
rect 504186 301258 504422 301494
rect 503866 300938 504102 301174
rect 504186 300938 504422 301174
rect 503866 267258 504102 267494
rect 504186 267258 504422 267494
rect 503866 266938 504102 267174
rect 504186 266938 504422 267174
rect 503866 233258 504102 233494
rect 504186 233258 504422 233494
rect 503866 232938 504102 233174
rect 504186 232938 504422 233174
rect 503866 199258 504102 199494
rect 504186 199258 504422 199494
rect 503866 198938 504102 199174
rect 504186 198938 504422 199174
rect 503866 165258 504102 165494
rect 504186 165258 504422 165494
rect 503866 164938 504102 165174
rect 504186 164938 504422 165174
rect 503866 131258 504102 131494
rect 504186 131258 504422 131494
rect 503866 130938 504102 131174
rect 504186 130938 504422 131174
rect 503866 97258 504102 97494
rect 504186 97258 504422 97494
rect 503866 96938 504102 97174
rect 504186 96938 504422 97174
rect 503866 63258 504102 63494
rect 504186 63258 504422 63494
rect 503866 62938 504102 63174
rect 504186 62938 504422 63174
rect 503866 29258 504102 29494
rect 504186 29258 504422 29494
rect 503866 28938 504102 29174
rect 504186 28938 504422 29174
rect 503866 -7302 504102 -7066
rect 504186 -7302 504422 -7066
rect 503866 -7622 504102 -7386
rect 504186 -7622 504422 -7386
rect 511826 704602 512062 704838
rect 512146 704602 512382 704838
rect 511826 704282 512062 704518
rect 512146 704282 512382 704518
rect 511826 683218 512062 683454
rect 512146 683218 512382 683454
rect 511826 682898 512062 683134
rect 512146 682898 512382 683134
rect 511826 649218 512062 649454
rect 512146 649218 512382 649454
rect 511826 648898 512062 649134
rect 512146 648898 512382 649134
rect 511826 615218 512062 615454
rect 512146 615218 512382 615454
rect 511826 614898 512062 615134
rect 512146 614898 512382 615134
rect 511826 581218 512062 581454
rect 512146 581218 512382 581454
rect 511826 580898 512062 581134
rect 512146 580898 512382 581134
rect 511826 547218 512062 547454
rect 512146 547218 512382 547454
rect 511826 546898 512062 547134
rect 512146 546898 512382 547134
rect 511826 513218 512062 513454
rect 512146 513218 512382 513454
rect 511826 512898 512062 513134
rect 512146 512898 512382 513134
rect 511826 479218 512062 479454
rect 512146 479218 512382 479454
rect 511826 478898 512062 479134
rect 512146 478898 512382 479134
rect 511826 445218 512062 445454
rect 512146 445218 512382 445454
rect 511826 444898 512062 445134
rect 512146 444898 512382 445134
rect 511826 411218 512062 411454
rect 512146 411218 512382 411454
rect 511826 410898 512062 411134
rect 512146 410898 512382 411134
rect 511826 377218 512062 377454
rect 512146 377218 512382 377454
rect 511826 376898 512062 377134
rect 512146 376898 512382 377134
rect 511826 343218 512062 343454
rect 512146 343218 512382 343454
rect 511826 342898 512062 343134
rect 512146 342898 512382 343134
rect 511826 309218 512062 309454
rect 512146 309218 512382 309454
rect 511826 308898 512062 309134
rect 512146 308898 512382 309134
rect 511826 275218 512062 275454
rect 512146 275218 512382 275454
rect 511826 274898 512062 275134
rect 512146 274898 512382 275134
rect 511826 241218 512062 241454
rect 512146 241218 512382 241454
rect 511826 240898 512062 241134
rect 512146 240898 512382 241134
rect 511826 207218 512062 207454
rect 512146 207218 512382 207454
rect 511826 206898 512062 207134
rect 512146 206898 512382 207134
rect 511826 173218 512062 173454
rect 512146 173218 512382 173454
rect 511826 172898 512062 173134
rect 512146 172898 512382 173134
rect 511826 139218 512062 139454
rect 512146 139218 512382 139454
rect 511826 138898 512062 139134
rect 512146 138898 512382 139134
rect 511826 105218 512062 105454
rect 512146 105218 512382 105454
rect 511826 104898 512062 105134
rect 512146 104898 512382 105134
rect 511826 71218 512062 71454
rect 512146 71218 512382 71454
rect 511826 70898 512062 71134
rect 512146 70898 512382 71134
rect 511826 37218 512062 37454
rect 512146 37218 512382 37454
rect 511826 36898 512062 37134
rect 512146 36898 512382 37134
rect 511826 3218 512062 3454
rect 512146 3218 512382 3454
rect 511826 2898 512062 3134
rect 512146 2898 512382 3134
rect 511826 -582 512062 -346
rect 512146 -582 512382 -346
rect 511826 -902 512062 -666
rect 512146 -902 512382 -666
rect 515546 705562 515782 705798
rect 515866 705562 516102 705798
rect 515546 705242 515782 705478
rect 515866 705242 516102 705478
rect 515546 686938 515782 687174
rect 515866 686938 516102 687174
rect 515546 686618 515782 686854
rect 515866 686618 516102 686854
rect 515546 652938 515782 653174
rect 515866 652938 516102 653174
rect 515546 652618 515782 652854
rect 515866 652618 516102 652854
rect 515546 618938 515782 619174
rect 515866 618938 516102 619174
rect 515546 618618 515782 618854
rect 515866 618618 516102 618854
rect 515546 584938 515782 585174
rect 515866 584938 516102 585174
rect 515546 584618 515782 584854
rect 515866 584618 516102 584854
rect 515546 550938 515782 551174
rect 515866 550938 516102 551174
rect 515546 550618 515782 550854
rect 515866 550618 516102 550854
rect 515546 516938 515782 517174
rect 515866 516938 516102 517174
rect 515546 516618 515782 516854
rect 515866 516618 516102 516854
rect 515546 482938 515782 483174
rect 515866 482938 516102 483174
rect 515546 482618 515782 482854
rect 515866 482618 516102 482854
rect 515546 448938 515782 449174
rect 515866 448938 516102 449174
rect 515546 448618 515782 448854
rect 515866 448618 516102 448854
rect 515546 414938 515782 415174
rect 515866 414938 516102 415174
rect 515546 414618 515782 414854
rect 515866 414618 516102 414854
rect 515546 380938 515782 381174
rect 515866 380938 516102 381174
rect 515546 380618 515782 380854
rect 515866 380618 516102 380854
rect 515546 346938 515782 347174
rect 515866 346938 516102 347174
rect 515546 346618 515782 346854
rect 515866 346618 516102 346854
rect 515546 312938 515782 313174
rect 515866 312938 516102 313174
rect 515546 312618 515782 312854
rect 515866 312618 516102 312854
rect 515546 278938 515782 279174
rect 515866 278938 516102 279174
rect 515546 278618 515782 278854
rect 515866 278618 516102 278854
rect 515546 244938 515782 245174
rect 515866 244938 516102 245174
rect 515546 244618 515782 244854
rect 515866 244618 516102 244854
rect 515546 210938 515782 211174
rect 515866 210938 516102 211174
rect 515546 210618 515782 210854
rect 515866 210618 516102 210854
rect 515546 176938 515782 177174
rect 515866 176938 516102 177174
rect 515546 176618 515782 176854
rect 515866 176618 516102 176854
rect 515546 142938 515782 143174
rect 515866 142938 516102 143174
rect 515546 142618 515782 142854
rect 515866 142618 516102 142854
rect 515546 108938 515782 109174
rect 515866 108938 516102 109174
rect 515546 108618 515782 108854
rect 515866 108618 516102 108854
rect 515546 74938 515782 75174
rect 515866 74938 516102 75174
rect 515546 74618 515782 74854
rect 515866 74618 516102 74854
rect 515546 40938 515782 41174
rect 515866 40938 516102 41174
rect 515546 40618 515782 40854
rect 515866 40618 516102 40854
rect 515546 6938 515782 7174
rect 515866 6938 516102 7174
rect 515546 6618 515782 6854
rect 515866 6618 516102 6854
rect 515546 -1542 515782 -1306
rect 515866 -1542 516102 -1306
rect 515546 -1862 515782 -1626
rect 515866 -1862 516102 -1626
rect 519266 706522 519502 706758
rect 519586 706522 519822 706758
rect 519266 706202 519502 706438
rect 519586 706202 519822 706438
rect 519266 690658 519502 690894
rect 519586 690658 519822 690894
rect 519266 690338 519502 690574
rect 519586 690338 519822 690574
rect 519266 656658 519502 656894
rect 519586 656658 519822 656894
rect 519266 656338 519502 656574
rect 519586 656338 519822 656574
rect 519266 622658 519502 622894
rect 519586 622658 519822 622894
rect 519266 622338 519502 622574
rect 519586 622338 519822 622574
rect 519266 588658 519502 588894
rect 519586 588658 519822 588894
rect 519266 588338 519502 588574
rect 519586 588338 519822 588574
rect 519266 554658 519502 554894
rect 519586 554658 519822 554894
rect 519266 554338 519502 554574
rect 519586 554338 519822 554574
rect 519266 520658 519502 520894
rect 519586 520658 519822 520894
rect 519266 520338 519502 520574
rect 519586 520338 519822 520574
rect 519266 486658 519502 486894
rect 519586 486658 519822 486894
rect 519266 486338 519502 486574
rect 519586 486338 519822 486574
rect 519266 452658 519502 452894
rect 519586 452658 519822 452894
rect 519266 452338 519502 452574
rect 519586 452338 519822 452574
rect 519266 418658 519502 418894
rect 519586 418658 519822 418894
rect 519266 418338 519502 418574
rect 519586 418338 519822 418574
rect 519266 384658 519502 384894
rect 519586 384658 519822 384894
rect 519266 384338 519502 384574
rect 519586 384338 519822 384574
rect 519266 350658 519502 350894
rect 519586 350658 519822 350894
rect 519266 350338 519502 350574
rect 519586 350338 519822 350574
rect 519266 316658 519502 316894
rect 519586 316658 519822 316894
rect 519266 316338 519502 316574
rect 519586 316338 519822 316574
rect 519266 282658 519502 282894
rect 519586 282658 519822 282894
rect 519266 282338 519502 282574
rect 519586 282338 519822 282574
rect 519266 248658 519502 248894
rect 519586 248658 519822 248894
rect 519266 248338 519502 248574
rect 519586 248338 519822 248574
rect 519266 214658 519502 214894
rect 519586 214658 519822 214894
rect 519266 214338 519502 214574
rect 519586 214338 519822 214574
rect 519266 180658 519502 180894
rect 519586 180658 519822 180894
rect 519266 180338 519502 180574
rect 519586 180338 519822 180574
rect 519266 146658 519502 146894
rect 519586 146658 519822 146894
rect 519266 146338 519502 146574
rect 519586 146338 519822 146574
rect 519266 112658 519502 112894
rect 519586 112658 519822 112894
rect 519266 112338 519502 112574
rect 519586 112338 519822 112574
rect 519266 78658 519502 78894
rect 519586 78658 519822 78894
rect 519266 78338 519502 78574
rect 519586 78338 519822 78574
rect 519266 44658 519502 44894
rect 519586 44658 519822 44894
rect 519266 44338 519502 44574
rect 519586 44338 519822 44574
rect 519266 10658 519502 10894
rect 519586 10658 519822 10894
rect 519266 10338 519502 10574
rect 519586 10338 519822 10574
rect 519266 -2502 519502 -2266
rect 519586 -2502 519822 -2266
rect 519266 -2822 519502 -2586
rect 519586 -2822 519822 -2586
rect 522986 707482 523222 707718
rect 523306 707482 523542 707718
rect 522986 707162 523222 707398
rect 523306 707162 523542 707398
rect 522986 694378 523222 694614
rect 523306 694378 523542 694614
rect 522986 694058 523222 694294
rect 523306 694058 523542 694294
rect 522986 660378 523222 660614
rect 523306 660378 523542 660614
rect 522986 660058 523222 660294
rect 523306 660058 523542 660294
rect 522986 626378 523222 626614
rect 523306 626378 523542 626614
rect 522986 626058 523222 626294
rect 523306 626058 523542 626294
rect 522986 592378 523222 592614
rect 523306 592378 523542 592614
rect 522986 592058 523222 592294
rect 523306 592058 523542 592294
rect 522986 558378 523222 558614
rect 523306 558378 523542 558614
rect 522986 558058 523222 558294
rect 523306 558058 523542 558294
rect 522986 524378 523222 524614
rect 523306 524378 523542 524614
rect 522986 524058 523222 524294
rect 523306 524058 523542 524294
rect 522986 490378 523222 490614
rect 523306 490378 523542 490614
rect 522986 490058 523222 490294
rect 523306 490058 523542 490294
rect 522986 456378 523222 456614
rect 523306 456378 523542 456614
rect 522986 456058 523222 456294
rect 523306 456058 523542 456294
rect 522986 422378 523222 422614
rect 523306 422378 523542 422614
rect 522986 422058 523222 422294
rect 523306 422058 523542 422294
rect 522986 388378 523222 388614
rect 523306 388378 523542 388614
rect 522986 388058 523222 388294
rect 523306 388058 523542 388294
rect 522986 354378 523222 354614
rect 523306 354378 523542 354614
rect 522986 354058 523222 354294
rect 523306 354058 523542 354294
rect 522986 320378 523222 320614
rect 523306 320378 523542 320614
rect 522986 320058 523222 320294
rect 523306 320058 523542 320294
rect 522986 286378 523222 286614
rect 523306 286378 523542 286614
rect 522986 286058 523222 286294
rect 523306 286058 523542 286294
rect 522986 252378 523222 252614
rect 523306 252378 523542 252614
rect 522986 252058 523222 252294
rect 523306 252058 523542 252294
rect 522986 218378 523222 218614
rect 523306 218378 523542 218614
rect 522986 218058 523222 218294
rect 523306 218058 523542 218294
rect 522986 184378 523222 184614
rect 523306 184378 523542 184614
rect 522986 184058 523222 184294
rect 523306 184058 523542 184294
rect 522986 150378 523222 150614
rect 523306 150378 523542 150614
rect 522986 150058 523222 150294
rect 523306 150058 523542 150294
rect 522986 116378 523222 116614
rect 523306 116378 523542 116614
rect 522986 116058 523222 116294
rect 523306 116058 523542 116294
rect 522986 82378 523222 82614
rect 523306 82378 523542 82614
rect 522986 82058 523222 82294
rect 523306 82058 523542 82294
rect 522986 48378 523222 48614
rect 523306 48378 523542 48614
rect 522986 48058 523222 48294
rect 523306 48058 523542 48294
rect 522986 14378 523222 14614
rect 523306 14378 523542 14614
rect 522986 14058 523222 14294
rect 523306 14058 523542 14294
rect 522986 -3462 523222 -3226
rect 523306 -3462 523542 -3226
rect 522986 -3782 523222 -3546
rect 523306 -3782 523542 -3546
rect 526706 708442 526942 708678
rect 527026 708442 527262 708678
rect 526706 708122 526942 708358
rect 527026 708122 527262 708358
rect 526706 698098 526942 698334
rect 527026 698098 527262 698334
rect 526706 697778 526942 698014
rect 527026 697778 527262 698014
rect 526706 664098 526942 664334
rect 527026 664098 527262 664334
rect 526706 663778 526942 664014
rect 527026 663778 527262 664014
rect 526706 630098 526942 630334
rect 527026 630098 527262 630334
rect 526706 629778 526942 630014
rect 527026 629778 527262 630014
rect 526706 596098 526942 596334
rect 527026 596098 527262 596334
rect 526706 595778 526942 596014
rect 527026 595778 527262 596014
rect 526706 562098 526942 562334
rect 527026 562098 527262 562334
rect 526706 561778 526942 562014
rect 527026 561778 527262 562014
rect 526706 528098 526942 528334
rect 527026 528098 527262 528334
rect 526706 527778 526942 528014
rect 527026 527778 527262 528014
rect 526706 494098 526942 494334
rect 527026 494098 527262 494334
rect 526706 493778 526942 494014
rect 527026 493778 527262 494014
rect 526706 460098 526942 460334
rect 527026 460098 527262 460334
rect 526706 459778 526942 460014
rect 527026 459778 527262 460014
rect 526706 426098 526942 426334
rect 527026 426098 527262 426334
rect 526706 425778 526942 426014
rect 527026 425778 527262 426014
rect 526706 392098 526942 392334
rect 527026 392098 527262 392334
rect 526706 391778 526942 392014
rect 527026 391778 527262 392014
rect 526706 358098 526942 358334
rect 527026 358098 527262 358334
rect 526706 357778 526942 358014
rect 527026 357778 527262 358014
rect 526706 324098 526942 324334
rect 527026 324098 527262 324334
rect 526706 323778 526942 324014
rect 527026 323778 527262 324014
rect 526706 290098 526942 290334
rect 527026 290098 527262 290334
rect 526706 289778 526942 290014
rect 527026 289778 527262 290014
rect 526706 256098 526942 256334
rect 527026 256098 527262 256334
rect 526706 255778 526942 256014
rect 527026 255778 527262 256014
rect 526706 222098 526942 222334
rect 527026 222098 527262 222334
rect 526706 221778 526942 222014
rect 527026 221778 527262 222014
rect 526706 188098 526942 188334
rect 527026 188098 527262 188334
rect 526706 187778 526942 188014
rect 527026 187778 527262 188014
rect 526706 154098 526942 154334
rect 527026 154098 527262 154334
rect 526706 153778 526942 154014
rect 527026 153778 527262 154014
rect 526706 120098 526942 120334
rect 527026 120098 527262 120334
rect 526706 119778 526942 120014
rect 527026 119778 527262 120014
rect 526706 86098 526942 86334
rect 527026 86098 527262 86334
rect 526706 85778 526942 86014
rect 527026 85778 527262 86014
rect 526706 52098 526942 52334
rect 527026 52098 527262 52334
rect 526706 51778 526942 52014
rect 527026 51778 527262 52014
rect 526706 18098 526942 18334
rect 527026 18098 527262 18334
rect 526706 17778 526942 18014
rect 527026 17778 527262 18014
rect 526706 -4422 526942 -4186
rect 527026 -4422 527262 -4186
rect 526706 -4742 526942 -4506
rect 527026 -4742 527262 -4506
rect 530426 709402 530662 709638
rect 530746 709402 530982 709638
rect 530426 709082 530662 709318
rect 530746 709082 530982 709318
rect 530426 667818 530662 668054
rect 530746 667818 530982 668054
rect 530426 667498 530662 667734
rect 530746 667498 530982 667734
rect 530426 633818 530662 634054
rect 530746 633818 530982 634054
rect 530426 633498 530662 633734
rect 530746 633498 530982 633734
rect 530426 599818 530662 600054
rect 530746 599818 530982 600054
rect 530426 599498 530662 599734
rect 530746 599498 530982 599734
rect 530426 565818 530662 566054
rect 530746 565818 530982 566054
rect 530426 565498 530662 565734
rect 530746 565498 530982 565734
rect 530426 531818 530662 532054
rect 530746 531818 530982 532054
rect 530426 531498 530662 531734
rect 530746 531498 530982 531734
rect 530426 497818 530662 498054
rect 530746 497818 530982 498054
rect 530426 497498 530662 497734
rect 530746 497498 530982 497734
rect 530426 463818 530662 464054
rect 530746 463818 530982 464054
rect 530426 463498 530662 463734
rect 530746 463498 530982 463734
rect 530426 429818 530662 430054
rect 530746 429818 530982 430054
rect 530426 429498 530662 429734
rect 530746 429498 530982 429734
rect 530426 395818 530662 396054
rect 530746 395818 530982 396054
rect 530426 395498 530662 395734
rect 530746 395498 530982 395734
rect 530426 361818 530662 362054
rect 530746 361818 530982 362054
rect 530426 361498 530662 361734
rect 530746 361498 530982 361734
rect 530426 327818 530662 328054
rect 530746 327818 530982 328054
rect 530426 327498 530662 327734
rect 530746 327498 530982 327734
rect 530426 293818 530662 294054
rect 530746 293818 530982 294054
rect 530426 293498 530662 293734
rect 530746 293498 530982 293734
rect 530426 259818 530662 260054
rect 530746 259818 530982 260054
rect 530426 259498 530662 259734
rect 530746 259498 530982 259734
rect 530426 225818 530662 226054
rect 530746 225818 530982 226054
rect 530426 225498 530662 225734
rect 530746 225498 530982 225734
rect 530426 191818 530662 192054
rect 530746 191818 530982 192054
rect 530426 191498 530662 191734
rect 530746 191498 530982 191734
rect 530426 157818 530662 158054
rect 530746 157818 530982 158054
rect 530426 157498 530662 157734
rect 530746 157498 530982 157734
rect 530426 123818 530662 124054
rect 530746 123818 530982 124054
rect 530426 123498 530662 123734
rect 530746 123498 530982 123734
rect 530426 89818 530662 90054
rect 530746 89818 530982 90054
rect 530426 89498 530662 89734
rect 530746 89498 530982 89734
rect 530426 55818 530662 56054
rect 530746 55818 530982 56054
rect 530426 55498 530662 55734
rect 530746 55498 530982 55734
rect 530426 21818 530662 22054
rect 530746 21818 530982 22054
rect 530426 21498 530662 21734
rect 530746 21498 530982 21734
rect 530426 -5382 530662 -5146
rect 530746 -5382 530982 -5146
rect 530426 -5702 530662 -5466
rect 530746 -5702 530982 -5466
rect 534146 710362 534382 710598
rect 534466 710362 534702 710598
rect 534146 710042 534382 710278
rect 534466 710042 534702 710278
rect 534146 671538 534382 671774
rect 534466 671538 534702 671774
rect 534146 671218 534382 671454
rect 534466 671218 534702 671454
rect 534146 637538 534382 637774
rect 534466 637538 534702 637774
rect 534146 637218 534382 637454
rect 534466 637218 534702 637454
rect 534146 603538 534382 603774
rect 534466 603538 534702 603774
rect 534146 603218 534382 603454
rect 534466 603218 534702 603454
rect 534146 569538 534382 569774
rect 534466 569538 534702 569774
rect 534146 569218 534382 569454
rect 534466 569218 534702 569454
rect 534146 535538 534382 535774
rect 534466 535538 534702 535774
rect 534146 535218 534382 535454
rect 534466 535218 534702 535454
rect 534146 501538 534382 501774
rect 534466 501538 534702 501774
rect 534146 501218 534382 501454
rect 534466 501218 534702 501454
rect 534146 467538 534382 467774
rect 534466 467538 534702 467774
rect 534146 467218 534382 467454
rect 534466 467218 534702 467454
rect 534146 433538 534382 433774
rect 534466 433538 534702 433774
rect 534146 433218 534382 433454
rect 534466 433218 534702 433454
rect 534146 399538 534382 399774
rect 534466 399538 534702 399774
rect 534146 399218 534382 399454
rect 534466 399218 534702 399454
rect 534146 365538 534382 365774
rect 534466 365538 534702 365774
rect 534146 365218 534382 365454
rect 534466 365218 534702 365454
rect 534146 331538 534382 331774
rect 534466 331538 534702 331774
rect 534146 331218 534382 331454
rect 534466 331218 534702 331454
rect 534146 297538 534382 297774
rect 534466 297538 534702 297774
rect 534146 297218 534382 297454
rect 534466 297218 534702 297454
rect 534146 263538 534382 263774
rect 534466 263538 534702 263774
rect 534146 263218 534382 263454
rect 534466 263218 534702 263454
rect 534146 229538 534382 229774
rect 534466 229538 534702 229774
rect 534146 229218 534382 229454
rect 534466 229218 534702 229454
rect 534146 195538 534382 195774
rect 534466 195538 534702 195774
rect 534146 195218 534382 195454
rect 534466 195218 534702 195454
rect 534146 161538 534382 161774
rect 534466 161538 534702 161774
rect 534146 161218 534382 161454
rect 534466 161218 534702 161454
rect 534146 127538 534382 127774
rect 534466 127538 534702 127774
rect 534146 127218 534382 127454
rect 534466 127218 534702 127454
rect 534146 93538 534382 93774
rect 534466 93538 534702 93774
rect 534146 93218 534382 93454
rect 534466 93218 534702 93454
rect 534146 59538 534382 59774
rect 534466 59538 534702 59774
rect 534146 59218 534382 59454
rect 534466 59218 534702 59454
rect 534146 25538 534382 25774
rect 534466 25538 534702 25774
rect 534146 25218 534382 25454
rect 534466 25218 534702 25454
rect 534146 -6342 534382 -6106
rect 534466 -6342 534702 -6106
rect 534146 -6662 534382 -6426
rect 534466 -6662 534702 -6426
rect 537866 711322 538102 711558
rect 538186 711322 538422 711558
rect 537866 711002 538102 711238
rect 538186 711002 538422 711238
rect 537866 675258 538102 675494
rect 538186 675258 538422 675494
rect 537866 674938 538102 675174
rect 538186 674938 538422 675174
rect 537866 641258 538102 641494
rect 538186 641258 538422 641494
rect 537866 640938 538102 641174
rect 538186 640938 538422 641174
rect 537866 607258 538102 607494
rect 538186 607258 538422 607494
rect 537866 606938 538102 607174
rect 538186 606938 538422 607174
rect 537866 573258 538102 573494
rect 538186 573258 538422 573494
rect 537866 572938 538102 573174
rect 538186 572938 538422 573174
rect 537866 539258 538102 539494
rect 538186 539258 538422 539494
rect 537866 538938 538102 539174
rect 538186 538938 538422 539174
rect 537866 505258 538102 505494
rect 538186 505258 538422 505494
rect 537866 504938 538102 505174
rect 538186 504938 538422 505174
rect 537866 471258 538102 471494
rect 538186 471258 538422 471494
rect 537866 470938 538102 471174
rect 538186 470938 538422 471174
rect 537866 437258 538102 437494
rect 538186 437258 538422 437494
rect 537866 436938 538102 437174
rect 538186 436938 538422 437174
rect 537866 403258 538102 403494
rect 538186 403258 538422 403494
rect 537866 402938 538102 403174
rect 538186 402938 538422 403174
rect 537866 369258 538102 369494
rect 538186 369258 538422 369494
rect 537866 368938 538102 369174
rect 538186 368938 538422 369174
rect 537866 335258 538102 335494
rect 538186 335258 538422 335494
rect 537866 334938 538102 335174
rect 538186 334938 538422 335174
rect 537866 301258 538102 301494
rect 538186 301258 538422 301494
rect 537866 300938 538102 301174
rect 538186 300938 538422 301174
rect 537866 267258 538102 267494
rect 538186 267258 538422 267494
rect 537866 266938 538102 267174
rect 538186 266938 538422 267174
rect 537866 233258 538102 233494
rect 538186 233258 538422 233494
rect 537866 232938 538102 233174
rect 538186 232938 538422 233174
rect 537866 199258 538102 199494
rect 538186 199258 538422 199494
rect 537866 198938 538102 199174
rect 538186 198938 538422 199174
rect 537866 165258 538102 165494
rect 538186 165258 538422 165494
rect 537866 164938 538102 165174
rect 538186 164938 538422 165174
rect 537866 131258 538102 131494
rect 538186 131258 538422 131494
rect 537866 130938 538102 131174
rect 538186 130938 538422 131174
rect 537866 97258 538102 97494
rect 538186 97258 538422 97494
rect 537866 96938 538102 97174
rect 538186 96938 538422 97174
rect 537866 63258 538102 63494
rect 538186 63258 538422 63494
rect 537866 62938 538102 63174
rect 538186 62938 538422 63174
rect 537866 29258 538102 29494
rect 538186 29258 538422 29494
rect 537866 28938 538102 29174
rect 538186 28938 538422 29174
rect 537866 -7302 538102 -7066
rect 538186 -7302 538422 -7066
rect 537866 -7622 538102 -7386
rect 538186 -7622 538422 -7386
rect 545826 704602 546062 704838
rect 546146 704602 546382 704838
rect 545826 704282 546062 704518
rect 546146 704282 546382 704518
rect 545826 683218 546062 683454
rect 546146 683218 546382 683454
rect 545826 682898 546062 683134
rect 546146 682898 546382 683134
rect 545826 649218 546062 649454
rect 546146 649218 546382 649454
rect 545826 648898 546062 649134
rect 546146 648898 546382 649134
rect 545826 615218 546062 615454
rect 546146 615218 546382 615454
rect 545826 614898 546062 615134
rect 546146 614898 546382 615134
rect 545826 581218 546062 581454
rect 546146 581218 546382 581454
rect 545826 580898 546062 581134
rect 546146 580898 546382 581134
rect 545826 547218 546062 547454
rect 546146 547218 546382 547454
rect 545826 546898 546062 547134
rect 546146 546898 546382 547134
rect 545826 513218 546062 513454
rect 546146 513218 546382 513454
rect 545826 512898 546062 513134
rect 546146 512898 546382 513134
rect 545826 479218 546062 479454
rect 546146 479218 546382 479454
rect 545826 478898 546062 479134
rect 546146 478898 546382 479134
rect 545826 445218 546062 445454
rect 546146 445218 546382 445454
rect 545826 444898 546062 445134
rect 546146 444898 546382 445134
rect 545826 411218 546062 411454
rect 546146 411218 546382 411454
rect 545826 410898 546062 411134
rect 546146 410898 546382 411134
rect 545826 377218 546062 377454
rect 546146 377218 546382 377454
rect 545826 376898 546062 377134
rect 546146 376898 546382 377134
rect 545826 343218 546062 343454
rect 546146 343218 546382 343454
rect 545826 342898 546062 343134
rect 546146 342898 546382 343134
rect 545826 309218 546062 309454
rect 546146 309218 546382 309454
rect 545826 308898 546062 309134
rect 546146 308898 546382 309134
rect 545826 275218 546062 275454
rect 546146 275218 546382 275454
rect 545826 274898 546062 275134
rect 546146 274898 546382 275134
rect 545826 241218 546062 241454
rect 546146 241218 546382 241454
rect 545826 240898 546062 241134
rect 546146 240898 546382 241134
rect 545826 207218 546062 207454
rect 546146 207218 546382 207454
rect 545826 206898 546062 207134
rect 546146 206898 546382 207134
rect 545826 173218 546062 173454
rect 546146 173218 546382 173454
rect 545826 172898 546062 173134
rect 546146 172898 546382 173134
rect 545826 139218 546062 139454
rect 546146 139218 546382 139454
rect 545826 138898 546062 139134
rect 546146 138898 546382 139134
rect 545826 105218 546062 105454
rect 546146 105218 546382 105454
rect 545826 104898 546062 105134
rect 546146 104898 546382 105134
rect 545826 71218 546062 71454
rect 546146 71218 546382 71454
rect 545826 70898 546062 71134
rect 546146 70898 546382 71134
rect 545826 37218 546062 37454
rect 546146 37218 546382 37454
rect 545826 36898 546062 37134
rect 546146 36898 546382 37134
rect 545826 3218 546062 3454
rect 546146 3218 546382 3454
rect 545826 2898 546062 3134
rect 546146 2898 546382 3134
rect 545826 -582 546062 -346
rect 546146 -582 546382 -346
rect 545826 -902 546062 -666
rect 546146 -902 546382 -666
rect 549546 705562 549782 705798
rect 549866 705562 550102 705798
rect 549546 705242 549782 705478
rect 549866 705242 550102 705478
rect 549546 686938 549782 687174
rect 549866 686938 550102 687174
rect 549546 686618 549782 686854
rect 549866 686618 550102 686854
rect 549546 652938 549782 653174
rect 549866 652938 550102 653174
rect 549546 652618 549782 652854
rect 549866 652618 550102 652854
rect 549546 618938 549782 619174
rect 549866 618938 550102 619174
rect 549546 618618 549782 618854
rect 549866 618618 550102 618854
rect 549546 584938 549782 585174
rect 549866 584938 550102 585174
rect 549546 584618 549782 584854
rect 549866 584618 550102 584854
rect 549546 550938 549782 551174
rect 549866 550938 550102 551174
rect 549546 550618 549782 550854
rect 549866 550618 550102 550854
rect 549546 516938 549782 517174
rect 549866 516938 550102 517174
rect 549546 516618 549782 516854
rect 549866 516618 550102 516854
rect 549546 482938 549782 483174
rect 549866 482938 550102 483174
rect 549546 482618 549782 482854
rect 549866 482618 550102 482854
rect 549546 448938 549782 449174
rect 549866 448938 550102 449174
rect 549546 448618 549782 448854
rect 549866 448618 550102 448854
rect 549546 414938 549782 415174
rect 549866 414938 550102 415174
rect 549546 414618 549782 414854
rect 549866 414618 550102 414854
rect 549546 380938 549782 381174
rect 549866 380938 550102 381174
rect 549546 380618 549782 380854
rect 549866 380618 550102 380854
rect 549546 346938 549782 347174
rect 549866 346938 550102 347174
rect 549546 346618 549782 346854
rect 549866 346618 550102 346854
rect 549546 312938 549782 313174
rect 549866 312938 550102 313174
rect 549546 312618 549782 312854
rect 549866 312618 550102 312854
rect 549546 278938 549782 279174
rect 549866 278938 550102 279174
rect 549546 278618 549782 278854
rect 549866 278618 550102 278854
rect 549546 244938 549782 245174
rect 549866 244938 550102 245174
rect 549546 244618 549782 244854
rect 549866 244618 550102 244854
rect 549546 210938 549782 211174
rect 549866 210938 550102 211174
rect 549546 210618 549782 210854
rect 549866 210618 550102 210854
rect 549546 176938 549782 177174
rect 549866 176938 550102 177174
rect 549546 176618 549782 176854
rect 549866 176618 550102 176854
rect 549546 142938 549782 143174
rect 549866 142938 550102 143174
rect 549546 142618 549782 142854
rect 549866 142618 550102 142854
rect 549546 108938 549782 109174
rect 549866 108938 550102 109174
rect 549546 108618 549782 108854
rect 549866 108618 550102 108854
rect 549546 74938 549782 75174
rect 549866 74938 550102 75174
rect 549546 74618 549782 74854
rect 549866 74618 550102 74854
rect 549546 40938 549782 41174
rect 549866 40938 550102 41174
rect 549546 40618 549782 40854
rect 549866 40618 550102 40854
rect 549546 6938 549782 7174
rect 549866 6938 550102 7174
rect 549546 6618 549782 6854
rect 549866 6618 550102 6854
rect 549546 -1542 549782 -1306
rect 549866 -1542 550102 -1306
rect 549546 -1862 549782 -1626
rect 549866 -1862 550102 -1626
rect 553266 706522 553502 706758
rect 553586 706522 553822 706758
rect 553266 706202 553502 706438
rect 553586 706202 553822 706438
rect 553266 690658 553502 690894
rect 553586 690658 553822 690894
rect 553266 690338 553502 690574
rect 553586 690338 553822 690574
rect 553266 656658 553502 656894
rect 553586 656658 553822 656894
rect 553266 656338 553502 656574
rect 553586 656338 553822 656574
rect 553266 622658 553502 622894
rect 553586 622658 553822 622894
rect 553266 622338 553502 622574
rect 553586 622338 553822 622574
rect 553266 588658 553502 588894
rect 553586 588658 553822 588894
rect 553266 588338 553502 588574
rect 553586 588338 553822 588574
rect 553266 554658 553502 554894
rect 553586 554658 553822 554894
rect 553266 554338 553502 554574
rect 553586 554338 553822 554574
rect 553266 520658 553502 520894
rect 553586 520658 553822 520894
rect 553266 520338 553502 520574
rect 553586 520338 553822 520574
rect 553266 486658 553502 486894
rect 553586 486658 553822 486894
rect 553266 486338 553502 486574
rect 553586 486338 553822 486574
rect 553266 452658 553502 452894
rect 553586 452658 553822 452894
rect 553266 452338 553502 452574
rect 553586 452338 553822 452574
rect 553266 418658 553502 418894
rect 553586 418658 553822 418894
rect 553266 418338 553502 418574
rect 553586 418338 553822 418574
rect 553266 384658 553502 384894
rect 553586 384658 553822 384894
rect 553266 384338 553502 384574
rect 553586 384338 553822 384574
rect 553266 350658 553502 350894
rect 553586 350658 553822 350894
rect 553266 350338 553502 350574
rect 553586 350338 553822 350574
rect 553266 316658 553502 316894
rect 553586 316658 553822 316894
rect 553266 316338 553502 316574
rect 553586 316338 553822 316574
rect 553266 282658 553502 282894
rect 553586 282658 553822 282894
rect 553266 282338 553502 282574
rect 553586 282338 553822 282574
rect 553266 248658 553502 248894
rect 553586 248658 553822 248894
rect 553266 248338 553502 248574
rect 553586 248338 553822 248574
rect 553266 214658 553502 214894
rect 553586 214658 553822 214894
rect 553266 214338 553502 214574
rect 553586 214338 553822 214574
rect 553266 180658 553502 180894
rect 553586 180658 553822 180894
rect 553266 180338 553502 180574
rect 553586 180338 553822 180574
rect 553266 146658 553502 146894
rect 553586 146658 553822 146894
rect 553266 146338 553502 146574
rect 553586 146338 553822 146574
rect 553266 112658 553502 112894
rect 553586 112658 553822 112894
rect 553266 112338 553502 112574
rect 553586 112338 553822 112574
rect 553266 78658 553502 78894
rect 553586 78658 553822 78894
rect 553266 78338 553502 78574
rect 553586 78338 553822 78574
rect 553266 44658 553502 44894
rect 553586 44658 553822 44894
rect 553266 44338 553502 44574
rect 553586 44338 553822 44574
rect 553266 10658 553502 10894
rect 553586 10658 553822 10894
rect 553266 10338 553502 10574
rect 553586 10338 553822 10574
rect 553266 -2502 553502 -2266
rect 553586 -2502 553822 -2266
rect 553266 -2822 553502 -2586
rect 553586 -2822 553822 -2586
rect 556986 707482 557222 707718
rect 557306 707482 557542 707718
rect 556986 707162 557222 707398
rect 557306 707162 557542 707398
rect 556986 694378 557222 694614
rect 557306 694378 557542 694614
rect 556986 694058 557222 694294
rect 557306 694058 557542 694294
rect 556986 660378 557222 660614
rect 557306 660378 557542 660614
rect 556986 660058 557222 660294
rect 557306 660058 557542 660294
rect 556986 626378 557222 626614
rect 557306 626378 557542 626614
rect 556986 626058 557222 626294
rect 557306 626058 557542 626294
rect 556986 592378 557222 592614
rect 557306 592378 557542 592614
rect 556986 592058 557222 592294
rect 557306 592058 557542 592294
rect 556986 558378 557222 558614
rect 557306 558378 557542 558614
rect 556986 558058 557222 558294
rect 557306 558058 557542 558294
rect 556986 524378 557222 524614
rect 557306 524378 557542 524614
rect 556986 524058 557222 524294
rect 557306 524058 557542 524294
rect 556986 490378 557222 490614
rect 557306 490378 557542 490614
rect 556986 490058 557222 490294
rect 557306 490058 557542 490294
rect 556986 456378 557222 456614
rect 557306 456378 557542 456614
rect 556986 456058 557222 456294
rect 557306 456058 557542 456294
rect 556986 422378 557222 422614
rect 557306 422378 557542 422614
rect 556986 422058 557222 422294
rect 557306 422058 557542 422294
rect 556986 388378 557222 388614
rect 557306 388378 557542 388614
rect 556986 388058 557222 388294
rect 557306 388058 557542 388294
rect 556986 354378 557222 354614
rect 557306 354378 557542 354614
rect 556986 354058 557222 354294
rect 557306 354058 557542 354294
rect 556986 320378 557222 320614
rect 557306 320378 557542 320614
rect 556986 320058 557222 320294
rect 557306 320058 557542 320294
rect 556986 286378 557222 286614
rect 557306 286378 557542 286614
rect 556986 286058 557222 286294
rect 557306 286058 557542 286294
rect 556986 252378 557222 252614
rect 557306 252378 557542 252614
rect 556986 252058 557222 252294
rect 557306 252058 557542 252294
rect 556986 218378 557222 218614
rect 557306 218378 557542 218614
rect 556986 218058 557222 218294
rect 557306 218058 557542 218294
rect 556986 184378 557222 184614
rect 557306 184378 557542 184614
rect 556986 184058 557222 184294
rect 557306 184058 557542 184294
rect 556986 150378 557222 150614
rect 557306 150378 557542 150614
rect 556986 150058 557222 150294
rect 557306 150058 557542 150294
rect 556986 116378 557222 116614
rect 557306 116378 557542 116614
rect 556986 116058 557222 116294
rect 557306 116058 557542 116294
rect 556986 82378 557222 82614
rect 557306 82378 557542 82614
rect 556986 82058 557222 82294
rect 557306 82058 557542 82294
rect 556986 48378 557222 48614
rect 557306 48378 557542 48614
rect 556986 48058 557222 48294
rect 557306 48058 557542 48294
rect 556986 14378 557222 14614
rect 557306 14378 557542 14614
rect 556986 14058 557222 14294
rect 557306 14058 557542 14294
rect 556986 -3462 557222 -3226
rect 557306 -3462 557542 -3226
rect 556986 -3782 557222 -3546
rect 557306 -3782 557542 -3546
rect 560706 708442 560942 708678
rect 561026 708442 561262 708678
rect 560706 708122 560942 708358
rect 561026 708122 561262 708358
rect 560706 698098 560942 698334
rect 561026 698098 561262 698334
rect 560706 697778 560942 698014
rect 561026 697778 561262 698014
rect 560706 664098 560942 664334
rect 561026 664098 561262 664334
rect 560706 663778 560942 664014
rect 561026 663778 561262 664014
rect 560706 630098 560942 630334
rect 561026 630098 561262 630334
rect 560706 629778 560942 630014
rect 561026 629778 561262 630014
rect 560706 596098 560942 596334
rect 561026 596098 561262 596334
rect 560706 595778 560942 596014
rect 561026 595778 561262 596014
rect 560706 562098 560942 562334
rect 561026 562098 561262 562334
rect 560706 561778 560942 562014
rect 561026 561778 561262 562014
rect 560706 528098 560942 528334
rect 561026 528098 561262 528334
rect 560706 527778 560942 528014
rect 561026 527778 561262 528014
rect 560706 494098 560942 494334
rect 561026 494098 561262 494334
rect 560706 493778 560942 494014
rect 561026 493778 561262 494014
rect 560706 460098 560942 460334
rect 561026 460098 561262 460334
rect 560706 459778 560942 460014
rect 561026 459778 561262 460014
rect 560706 426098 560942 426334
rect 561026 426098 561262 426334
rect 560706 425778 560942 426014
rect 561026 425778 561262 426014
rect 560706 392098 560942 392334
rect 561026 392098 561262 392334
rect 560706 391778 560942 392014
rect 561026 391778 561262 392014
rect 560706 358098 560942 358334
rect 561026 358098 561262 358334
rect 560706 357778 560942 358014
rect 561026 357778 561262 358014
rect 560706 324098 560942 324334
rect 561026 324098 561262 324334
rect 560706 323778 560942 324014
rect 561026 323778 561262 324014
rect 560706 290098 560942 290334
rect 561026 290098 561262 290334
rect 560706 289778 560942 290014
rect 561026 289778 561262 290014
rect 560706 256098 560942 256334
rect 561026 256098 561262 256334
rect 560706 255778 560942 256014
rect 561026 255778 561262 256014
rect 560706 222098 560942 222334
rect 561026 222098 561262 222334
rect 560706 221778 560942 222014
rect 561026 221778 561262 222014
rect 560706 188098 560942 188334
rect 561026 188098 561262 188334
rect 560706 187778 560942 188014
rect 561026 187778 561262 188014
rect 560706 154098 560942 154334
rect 561026 154098 561262 154334
rect 560706 153778 560942 154014
rect 561026 153778 561262 154014
rect 560706 120098 560942 120334
rect 561026 120098 561262 120334
rect 560706 119778 560942 120014
rect 561026 119778 561262 120014
rect 560706 86098 560942 86334
rect 561026 86098 561262 86334
rect 560706 85778 560942 86014
rect 561026 85778 561262 86014
rect 560706 52098 560942 52334
rect 561026 52098 561262 52334
rect 560706 51778 560942 52014
rect 561026 51778 561262 52014
rect 560706 18098 560942 18334
rect 561026 18098 561262 18334
rect 560706 17778 560942 18014
rect 561026 17778 561262 18014
rect 560706 -4422 560942 -4186
rect 561026 -4422 561262 -4186
rect 560706 -4742 560942 -4506
rect 561026 -4742 561262 -4506
rect 564426 709402 564662 709638
rect 564746 709402 564982 709638
rect 564426 709082 564662 709318
rect 564746 709082 564982 709318
rect 564426 667818 564662 668054
rect 564746 667818 564982 668054
rect 564426 667498 564662 667734
rect 564746 667498 564982 667734
rect 564426 633818 564662 634054
rect 564746 633818 564982 634054
rect 564426 633498 564662 633734
rect 564746 633498 564982 633734
rect 564426 599818 564662 600054
rect 564746 599818 564982 600054
rect 564426 599498 564662 599734
rect 564746 599498 564982 599734
rect 564426 565818 564662 566054
rect 564746 565818 564982 566054
rect 564426 565498 564662 565734
rect 564746 565498 564982 565734
rect 564426 531818 564662 532054
rect 564746 531818 564982 532054
rect 564426 531498 564662 531734
rect 564746 531498 564982 531734
rect 564426 497818 564662 498054
rect 564746 497818 564982 498054
rect 564426 497498 564662 497734
rect 564746 497498 564982 497734
rect 564426 463818 564662 464054
rect 564746 463818 564982 464054
rect 564426 463498 564662 463734
rect 564746 463498 564982 463734
rect 564426 429818 564662 430054
rect 564746 429818 564982 430054
rect 564426 429498 564662 429734
rect 564746 429498 564982 429734
rect 564426 395818 564662 396054
rect 564746 395818 564982 396054
rect 564426 395498 564662 395734
rect 564746 395498 564982 395734
rect 564426 361818 564662 362054
rect 564746 361818 564982 362054
rect 564426 361498 564662 361734
rect 564746 361498 564982 361734
rect 564426 327818 564662 328054
rect 564746 327818 564982 328054
rect 564426 327498 564662 327734
rect 564746 327498 564982 327734
rect 564426 293818 564662 294054
rect 564746 293818 564982 294054
rect 564426 293498 564662 293734
rect 564746 293498 564982 293734
rect 564426 259818 564662 260054
rect 564746 259818 564982 260054
rect 564426 259498 564662 259734
rect 564746 259498 564982 259734
rect 564426 225818 564662 226054
rect 564746 225818 564982 226054
rect 564426 225498 564662 225734
rect 564746 225498 564982 225734
rect 564426 191818 564662 192054
rect 564746 191818 564982 192054
rect 564426 191498 564662 191734
rect 564746 191498 564982 191734
rect 564426 157818 564662 158054
rect 564746 157818 564982 158054
rect 564426 157498 564662 157734
rect 564746 157498 564982 157734
rect 564426 123818 564662 124054
rect 564746 123818 564982 124054
rect 564426 123498 564662 123734
rect 564746 123498 564982 123734
rect 564426 89818 564662 90054
rect 564746 89818 564982 90054
rect 564426 89498 564662 89734
rect 564746 89498 564982 89734
rect 564426 55818 564662 56054
rect 564746 55818 564982 56054
rect 564426 55498 564662 55734
rect 564746 55498 564982 55734
rect 564426 21818 564662 22054
rect 564746 21818 564982 22054
rect 564426 21498 564662 21734
rect 564746 21498 564982 21734
rect 564426 -5382 564662 -5146
rect 564746 -5382 564982 -5146
rect 564426 -5702 564662 -5466
rect 564746 -5702 564982 -5466
rect 568146 710362 568382 710598
rect 568466 710362 568702 710598
rect 568146 710042 568382 710278
rect 568466 710042 568702 710278
rect 568146 671538 568382 671774
rect 568466 671538 568702 671774
rect 568146 671218 568382 671454
rect 568466 671218 568702 671454
rect 568146 637538 568382 637774
rect 568466 637538 568702 637774
rect 568146 637218 568382 637454
rect 568466 637218 568702 637454
rect 568146 603538 568382 603774
rect 568466 603538 568702 603774
rect 568146 603218 568382 603454
rect 568466 603218 568702 603454
rect 568146 569538 568382 569774
rect 568466 569538 568702 569774
rect 568146 569218 568382 569454
rect 568466 569218 568702 569454
rect 568146 535538 568382 535774
rect 568466 535538 568702 535774
rect 568146 535218 568382 535454
rect 568466 535218 568702 535454
rect 568146 501538 568382 501774
rect 568466 501538 568702 501774
rect 568146 501218 568382 501454
rect 568466 501218 568702 501454
rect 568146 467538 568382 467774
rect 568466 467538 568702 467774
rect 568146 467218 568382 467454
rect 568466 467218 568702 467454
rect 568146 433538 568382 433774
rect 568466 433538 568702 433774
rect 568146 433218 568382 433454
rect 568466 433218 568702 433454
rect 568146 399538 568382 399774
rect 568466 399538 568702 399774
rect 568146 399218 568382 399454
rect 568466 399218 568702 399454
rect 568146 365538 568382 365774
rect 568466 365538 568702 365774
rect 568146 365218 568382 365454
rect 568466 365218 568702 365454
rect 568146 331538 568382 331774
rect 568466 331538 568702 331774
rect 568146 331218 568382 331454
rect 568466 331218 568702 331454
rect 568146 297538 568382 297774
rect 568466 297538 568702 297774
rect 568146 297218 568382 297454
rect 568466 297218 568702 297454
rect 568146 263538 568382 263774
rect 568466 263538 568702 263774
rect 568146 263218 568382 263454
rect 568466 263218 568702 263454
rect 568146 229538 568382 229774
rect 568466 229538 568702 229774
rect 568146 229218 568382 229454
rect 568466 229218 568702 229454
rect 568146 195538 568382 195774
rect 568466 195538 568702 195774
rect 568146 195218 568382 195454
rect 568466 195218 568702 195454
rect 568146 161538 568382 161774
rect 568466 161538 568702 161774
rect 568146 161218 568382 161454
rect 568466 161218 568702 161454
rect 568146 127538 568382 127774
rect 568466 127538 568702 127774
rect 568146 127218 568382 127454
rect 568466 127218 568702 127454
rect 568146 93538 568382 93774
rect 568466 93538 568702 93774
rect 568146 93218 568382 93454
rect 568466 93218 568702 93454
rect 568146 59538 568382 59774
rect 568466 59538 568702 59774
rect 568146 59218 568382 59454
rect 568466 59218 568702 59454
rect 568146 25538 568382 25774
rect 568466 25538 568702 25774
rect 568146 25218 568382 25454
rect 568466 25218 568702 25454
rect 568146 -6342 568382 -6106
rect 568466 -6342 568702 -6106
rect 568146 -6662 568382 -6426
rect 568466 -6662 568702 -6426
rect 571866 711322 572102 711558
rect 572186 711322 572422 711558
rect 571866 711002 572102 711238
rect 572186 711002 572422 711238
rect 571866 675258 572102 675494
rect 572186 675258 572422 675494
rect 571866 674938 572102 675174
rect 572186 674938 572422 675174
rect 571866 641258 572102 641494
rect 572186 641258 572422 641494
rect 571866 640938 572102 641174
rect 572186 640938 572422 641174
rect 571866 607258 572102 607494
rect 572186 607258 572422 607494
rect 571866 606938 572102 607174
rect 572186 606938 572422 607174
rect 571866 573258 572102 573494
rect 572186 573258 572422 573494
rect 571866 572938 572102 573174
rect 572186 572938 572422 573174
rect 571866 539258 572102 539494
rect 572186 539258 572422 539494
rect 571866 538938 572102 539174
rect 572186 538938 572422 539174
rect 571866 505258 572102 505494
rect 572186 505258 572422 505494
rect 571866 504938 572102 505174
rect 572186 504938 572422 505174
rect 571866 471258 572102 471494
rect 572186 471258 572422 471494
rect 571866 470938 572102 471174
rect 572186 470938 572422 471174
rect 571866 437258 572102 437494
rect 572186 437258 572422 437494
rect 571866 436938 572102 437174
rect 572186 436938 572422 437174
rect 571866 403258 572102 403494
rect 572186 403258 572422 403494
rect 571866 402938 572102 403174
rect 572186 402938 572422 403174
rect 571866 369258 572102 369494
rect 572186 369258 572422 369494
rect 571866 368938 572102 369174
rect 572186 368938 572422 369174
rect 571866 335258 572102 335494
rect 572186 335258 572422 335494
rect 571866 334938 572102 335174
rect 572186 334938 572422 335174
rect 571866 301258 572102 301494
rect 572186 301258 572422 301494
rect 571866 300938 572102 301174
rect 572186 300938 572422 301174
rect 571866 267258 572102 267494
rect 572186 267258 572422 267494
rect 571866 266938 572102 267174
rect 572186 266938 572422 267174
rect 571866 233258 572102 233494
rect 572186 233258 572422 233494
rect 571866 232938 572102 233174
rect 572186 232938 572422 233174
rect 571866 199258 572102 199494
rect 572186 199258 572422 199494
rect 571866 198938 572102 199174
rect 572186 198938 572422 199174
rect 571866 165258 572102 165494
rect 572186 165258 572422 165494
rect 571866 164938 572102 165174
rect 572186 164938 572422 165174
rect 571866 131258 572102 131494
rect 572186 131258 572422 131494
rect 571866 130938 572102 131174
rect 572186 130938 572422 131174
rect 571866 97258 572102 97494
rect 572186 97258 572422 97494
rect 571866 96938 572102 97174
rect 572186 96938 572422 97174
rect 571866 63258 572102 63494
rect 572186 63258 572422 63494
rect 571866 62938 572102 63174
rect 572186 62938 572422 63174
rect 571866 29258 572102 29494
rect 572186 29258 572422 29494
rect 571866 28938 572102 29174
rect 572186 28938 572422 29174
rect 571866 -7302 572102 -7066
rect 572186 -7302 572422 -7066
rect 571866 -7622 572102 -7386
rect 572186 -7622 572422 -7386
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 579826 704602 580062 704838
rect 580146 704602 580382 704838
rect 579826 704282 580062 704518
rect 580146 704282 580382 704518
rect 579826 683218 580062 683454
rect 580146 683218 580382 683454
rect 579826 682898 580062 683134
rect 580146 682898 580382 683134
rect 579826 649218 580062 649454
rect 580146 649218 580382 649454
rect 579826 648898 580062 649134
rect 580146 648898 580382 649134
rect 579826 615218 580062 615454
rect 580146 615218 580382 615454
rect 579826 614898 580062 615134
rect 580146 614898 580382 615134
rect 579826 581218 580062 581454
rect 580146 581218 580382 581454
rect 579826 580898 580062 581134
rect 580146 580898 580382 581134
rect 579826 547218 580062 547454
rect 580146 547218 580382 547454
rect 579826 546898 580062 547134
rect 580146 546898 580382 547134
rect 579826 513218 580062 513454
rect 580146 513218 580382 513454
rect 579826 512898 580062 513134
rect 580146 512898 580382 513134
rect 579826 479218 580062 479454
rect 580146 479218 580382 479454
rect 579826 478898 580062 479134
rect 580146 478898 580382 479134
rect 579826 445218 580062 445454
rect 580146 445218 580382 445454
rect 579826 444898 580062 445134
rect 580146 444898 580382 445134
rect 579826 411218 580062 411454
rect 580146 411218 580382 411454
rect 579826 410898 580062 411134
rect 580146 410898 580382 411134
rect 579826 377218 580062 377454
rect 580146 377218 580382 377454
rect 579826 376898 580062 377134
rect 580146 376898 580382 377134
rect 579826 343218 580062 343454
rect 580146 343218 580382 343454
rect 579826 342898 580062 343134
rect 580146 342898 580382 343134
rect 579826 309218 580062 309454
rect 580146 309218 580382 309454
rect 579826 308898 580062 309134
rect 580146 308898 580382 309134
rect 579826 275218 580062 275454
rect 580146 275218 580382 275454
rect 579826 274898 580062 275134
rect 580146 274898 580382 275134
rect 579826 241218 580062 241454
rect 580146 241218 580382 241454
rect 579826 240898 580062 241134
rect 580146 240898 580382 241134
rect 579826 207218 580062 207454
rect 580146 207218 580382 207454
rect 579826 206898 580062 207134
rect 580146 206898 580382 207134
rect 579826 173218 580062 173454
rect 580146 173218 580382 173454
rect 579826 172898 580062 173134
rect 580146 172898 580382 173134
rect 579826 139218 580062 139454
rect 580146 139218 580382 139454
rect 579826 138898 580062 139134
rect 580146 138898 580382 139134
rect 579826 105218 580062 105454
rect 580146 105218 580382 105454
rect 579826 104898 580062 105134
rect 580146 104898 580382 105134
rect 579826 71218 580062 71454
rect 580146 71218 580382 71454
rect 579826 70898 580062 71134
rect 580146 70898 580382 71134
rect 579826 37218 580062 37454
rect 580146 37218 580382 37454
rect 579826 36898 580062 37134
rect 580146 36898 580382 37134
rect 579826 3218 580062 3454
rect 580146 3218 580382 3454
rect 579826 2898 580062 3134
rect 580146 2898 580382 3134
rect 579826 -582 580062 -346
rect 580146 -582 580382 -346
rect 579826 -902 580062 -666
rect 580146 -902 580382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 683218 585578 683454
rect 585662 683218 585898 683454
rect 585342 682898 585578 683134
rect 585662 682898 585898 683134
rect 585342 649218 585578 649454
rect 585662 649218 585898 649454
rect 585342 648898 585578 649134
rect 585662 648898 585898 649134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 581218 585578 581454
rect 585662 581218 585898 581454
rect 585342 580898 585578 581134
rect 585662 580898 585898 581134
rect 585342 547218 585578 547454
rect 585662 547218 585898 547454
rect 585342 546898 585578 547134
rect 585662 546898 585898 547134
rect 585342 513218 585578 513454
rect 585662 513218 585898 513454
rect 585342 512898 585578 513134
rect 585662 512898 585898 513134
rect 585342 479218 585578 479454
rect 585662 479218 585898 479454
rect 585342 478898 585578 479134
rect 585662 478898 585898 479134
rect 585342 445218 585578 445454
rect 585662 445218 585898 445454
rect 585342 444898 585578 445134
rect 585662 444898 585898 445134
rect 585342 411218 585578 411454
rect 585662 411218 585898 411454
rect 585342 410898 585578 411134
rect 585662 410898 585898 411134
rect 585342 377218 585578 377454
rect 585662 377218 585898 377454
rect 585342 376898 585578 377134
rect 585662 376898 585898 377134
rect 585342 343218 585578 343454
rect 585662 343218 585898 343454
rect 585342 342898 585578 343134
rect 585662 342898 585898 343134
rect 585342 309218 585578 309454
rect 585662 309218 585898 309454
rect 585342 308898 585578 309134
rect 585662 308898 585898 309134
rect 585342 275218 585578 275454
rect 585662 275218 585898 275454
rect 585342 274898 585578 275134
rect 585662 274898 585898 275134
rect 585342 241218 585578 241454
rect 585662 241218 585898 241454
rect 585342 240898 585578 241134
rect 585662 240898 585898 241134
rect 585342 207218 585578 207454
rect 585662 207218 585898 207454
rect 585342 206898 585578 207134
rect 585662 206898 585898 207134
rect 585342 173218 585578 173454
rect 585662 173218 585898 173454
rect 585342 172898 585578 173134
rect 585662 172898 585898 173134
rect 585342 139218 585578 139454
rect 585662 139218 585898 139454
rect 585342 138898 585578 139134
rect 585662 138898 585898 139134
rect 585342 105218 585578 105454
rect 585662 105218 585898 105454
rect 585342 104898 585578 105134
rect 585662 104898 585898 105134
rect 585342 71218 585578 71454
rect 585662 71218 585898 71454
rect 585342 70898 585578 71134
rect 585662 70898 585898 71134
rect 585342 37218 585578 37454
rect 585662 37218 585898 37454
rect 585342 36898 585578 37134
rect 585662 36898 585898 37134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 686938 586538 687174
rect 586622 686938 586858 687174
rect 586302 686618 586538 686854
rect 586622 686618 586858 686854
rect 586302 652938 586538 653174
rect 586622 652938 586858 653174
rect 586302 652618 586538 652854
rect 586622 652618 586858 652854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 584938 586538 585174
rect 586622 584938 586858 585174
rect 586302 584618 586538 584854
rect 586622 584618 586858 584854
rect 586302 550938 586538 551174
rect 586622 550938 586858 551174
rect 586302 550618 586538 550854
rect 586622 550618 586858 550854
rect 586302 516938 586538 517174
rect 586622 516938 586858 517174
rect 586302 516618 586538 516854
rect 586622 516618 586858 516854
rect 586302 482938 586538 483174
rect 586622 482938 586858 483174
rect 586302 482618 586538 482854
rect 586622 482618 586858 482854
rect 586302 448938 586538 449174
rect 586622 448938 586858 449174
rect 586302 448618 586538 448854
rect 586622 448618 586858 448854
rect 586302 414938 586538 415174
rect 586622 414938 586858 415174
rect 586302 414618 586538 414854
rect 586622 414618 586858 414854
rect 586302 380938 586538 381174
rect 586622 380938 586858 381174
rect 586302 380618 586538 380854
rect 586622 380618 586858 380854
rect 586302 346938 586538 347174
rect 586622 346938 586858 347174
rect 586302 346618 586538 346854
rect 586622 346618 586858 346854
rect 586302 312938 586538 313174
rect 586622 312938 586858 313174
rect 586302 312618 586538 312854
rect 586622 312618 586858 312854
rect 586302 278938 586538 279174
rect 586622 278938 586858 279174
rect 586302 278618 586538 278854
rect 586622 278618 586858 278854
rect 586302 244938 586538 245174
rect 586622 244938 586858 245174
rect 586302 244618 586538 244854
rect 586622 244618 586858 244854
rect 586302 210938 586538 211174
rect 586622 210938 586858 211174
rect 586302 210618 586538 210854
rect 586622 210618 586858 210854
rect 586302 176938 586538 177174
rect 586622 176938 586858 177174
rect 586302 176618 586538 176854
rect 586622 176618 586858 176854
rect 586302 142938 586538 143174
rect 586622 142938 586858 143174
rect 586302 142618 586538 142854
rect 586622 142618 586858 142854
rect 586302 108938 586538 109174
rect 586622 108938 586858 109174
rect 586302 108618 586538 108854
rect 586622 108618 586858 108854
rect 586302 74938 586538 75174
rect 586622 74938 586858 75174
rect 586302 74618 586538 74854
rect 586622 74618 586858 74854
rect 586302 40938 586538 41174
rect 586622 40938 586858 41174
rect 586302 40618 586538 40854
rect 586622 40618 586858 40854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690658 587498 690894
rect 587582 690658 587818 690894
rect 587262 690338 587498 690574
rect 587582 690338 587818 690574
rect 587262 656658 587498 656894
rect 587582 656658 587818 656894
rect 587262 656338 587498 656574
rect 587582 656338 587818 656574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 588658 587498 588894
rect 587582 588658 587818 588894
rect 587262 588338 587498 588574
rect 587582 588338 587818 588574
rect 587262 554658 587498 554894
rect 587582 554658 587818 554894
rect 587262 554338 587498 554574
rect 587582 554338 587818 554574
rect 587262 520658 587498 520894
rect 587582 520658 587818 520894
rect 587262 520338 587498 520574
rect 587582 520338 587818 520574
rect 587262 486658 587498 486894
rect 587582 486658 587818 486894
rect 587262 486338 587498 486574
rect 587582 486338 587818 486574
rect 587262 452658 587498 452894
rect 587582 452658 587818 452894
rect 587262 452338 587498 452574
rect 587582 452338 587818 452574
rect 587262 418658 587498 418894
rect 587582 418658 587818 418894
rect 587262 418338 587498 418574
rect 587582 418338 587818 418574
rect 587262 384658 587498 384894
rect 587582 384658 587818 384894
rect 587262 384338 587498 384574
rect 587582 384338 587818 384574
rect 587262 350658 587498 350894
rect 587582 350658 587818 350894
rect 587262 350338 587498 350574
rect 587582 350338 587818 350574
rect 587262 316658 587498 316894
rect 587582 316658 587818 316894
rect 587262 316338 587498 316574
rect 587582 316338 587818 316574
rect 587262 282658 587498 282894
rect 587582 282658 587818 282894
rect 587262 282338 587498 282574
rect 587582 282338 587818 282574
rect 587262 248658 587498 248894
rect 587582 248658 587818 248894
rect 587262 248338 587498 248574
rect 587582 248338 587818 248574
rect 587262 214658 587498 214894
rect 587582 214658 587818 214894
rect 587262 214338 587498 214574
rect 587582 214338 587818 214574
rect 587262 180658 587498 180894
rect 587582 180658 587818 180894
rect 587262 180338 587498 180574
rect 587582 180338 587818 180574
rect 587262 146658 587498 146894
rect 587582 146658 587818 146894
rect 587262 146338 587498 146574
rect 587582 146338 587818 146574
rect 587262 112658 587498 112894
rect 587582 112658 587818 112894
rect 587262 112338 587498 112574
rect 587582 112338 587818 112574
rect 587262 78658 587498 78894
rect 587582 78658 587818 78894
rect 587262 78338 587498 78574
rect 587582 78338 587818 78574
rect 587262 44658 587498 44894
rect 587582 44658 587818 44894
rect 587262 44338 587498 44574
rect 587582 44338 587818 44574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 694378 588458 694614
rect 588542 694378 588778 694614
rect 588222 694058 588458 694294
rect 588542 694058 588778 694294
rect 588222 660378 588458 660614
rect 588542 660378 588778 660614
rect 588222 660058 588458 660294
rect 588542 660058 588778 660294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 592378 588458 592614
rect 588542 592378 588778 592614
rect 588222 592058 588458 592294
rect 588542 592058 588778 592294
rect 588222 558378 588458 558614
rect 588542 558378 588778 558614
rect 588222 558058 588458 558294
rect 588542 558058 588778 558294
rect 588222 524378 588458 524614
rect 588542 524378 588778 524614
rect 588222 524058 588458 524294
rect 588542 524058 588778 524294
rect 588222 490378 588458 490614
rect 588542 490378 588778 490614
rect 588222 490058 588458 490294
rect 588542 490058 588778 490294
rect 588222 456378 588458 456614
rect 588542 456378 588778 456614
rect 588222 456058 588458 456294
rect 588542 456058 588778 456294
rect 588222 422378 588458 422614
rect 588542 422378 588778 422614
rect 588222 422058 588458 422294
rect 588542 422058 588778 422294
rect 588222 388378 588458 388614
rect 588542 388378 588778 388614
rect 588222 388058 588458 388294
rect 588542 388058 588778 388294
rect 588222 354378 588458 354614
rect 588542 354378 588778 354614
rect 588222 354058 588458 354294
rect 588542 354058 588778 354294
rect 588222 320378 588458 320614
rect 588542 320378 588778 320614
rect 588222 320058 588458 320294
rect 588542 320058 588778 320294
rect 588222 286378 588458 286614
rect 588542 286378 588778 286614
rect 588222 286058 588458 286294
rect 588542 286058 588778 286294
rect 588222 252378 588458 252614
rect 588542 252378 588778 252614
rect 588222 252058 588458 252294
rect 588542 252058 588778 252294
rect 588222 218378 588458 218614
rect 588542 218378 588778 218614
rect 588222 218058 588458 218294
rect 588542 218058 588778 218294
rect 588222 184378 588458 184614
rect 588542 184378 588778 184614
rect 588222 184058 588458 184294
rect 588542 184058 588778 184294
rect 588222 150378 588458 150614
rect 588542 150378 588778 150614
rect 588222 150058 588458 150294
rect 588542 150058 588778 150294
rect 588222 116378 588458 116614
rect 588542 116378 588778 116614
rect 588222 116058 588458 116294
rect 588542 116058 588778 116294
rect 588222 82378 588458 82614
rect 588542 82378 588778 82614
rect 588222 82058 588458 82294
rect 588542 82058 588778 82294
rect 588222 48378 588458 48614
rect 588542 48378 588778 48614
rect 588222 48058 588458 48294
rect 588542 48058 588778 48294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 698098 589418 698334
rect 589502 698098 589738 698334
rect 589182 697778 589418 698014
rect 589502 697778 589738 698014
rect 589182 664098 589418 664334
rect 589502 664098 589738 664334
rect 589182 663778 589418 664014
rect 589502 663778 589738 664014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 596098 589418 596334
rect 589502 596098 589738 596334
rect 589182 595778 589418 596014
rect 589502 595778 589738 596014
rect 589182 562098 589418 562334
rect 589502 562098 589738 562334
rect 589182 561778 589418 562014
rect 589502 561778 589738 562014
rect 589182 528098 589418 528334
rect 589502 528098 589738 528334
rect 589182 527778 589418 528014
rect 589502 527778 589738 528014
rect 589182 494098 589418 494334
rect 589502 494098 589738 494334
rect 589182 493778 589418 494014
rect 589502 493778 589738 494014
rect 589182 460098 589418 460334
rect 589502 460098 589738 460334
rect 589182 459778 589418 460014
rect 589502 459778 589738 460014
rect 589182 426098 589418 426334
rect 589502 426098 589738 426334
rect 589182 425778 589418 426014
rect 589502 425778 589738 426014
rect 589182 392098 589418 392334
rect 589502 392098 589738 392334
rect 589182 391778 589418 392014
rect 589502 391778 589738 392014
rect 589182 358098 589418 358334
rect 589502 358098 589738 358334
rect 589182 357778 589418 358014
rect 589502 357778 589738 358014
rect 589182 324098 589418 324334
rect 589502 324098 589738 324334
rect 589182 323778 589418 324014
rect 589502 323778 589738 324014
rect 589182 290098 589418 290334
rect 589502 290098 589738 290334
rect 589182 289778 589418 290014
rect 589502 289778 589738 290014
rect 589182 256098 589418 256334
rect 589502 256098 589738 256334
rect 589182 255778 589418 256014
rect 589502 255778 589738 256014
rect 589182 222098 589418 222334
rect 589502 222098 589738 222334
rect 589182 221778 589418 222014
rect 589502 221778 589738 222014
rect 589182 188098 589418 188334
rect 589502 188098 589738 188334
rect 589182 187778 589418 188014
rect 589502 187778 589738 188014
rect 589182 154098 589418 154334
rect 589502 154098 589738 154334
rect 589182 153778 589418 154014
rect 589502 153778 589738 154014
rect 589182 120098 589418 120334
rect 589502 120098 589738 120334
rect 589182 119778 589418 120014
rect 589502 119778 589738 120014
rect 589182 86098 589418 86334
rect 589502 86098 589738 86334
rect 589182 85778 589418 86014
rect 589502 85778 589738 86014
rect 589182 52098 589418 52334
rect 589502 52098 589738 52334
rect 589182 51778 589418 52014
rect 589502 51778 589738 52014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 667818 590378 668054
rect 590462 667818 590698 668054
rect 590142 667498 590378 667734
rect 590462 667498 590698 667734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 599818 590378 600054
rect 590462 599818 590698 600054
rect 590142 599498 590378 599734
rect 590462 599498 590698 599734
rect 590142 565818 590378 566054
rect 590462 565818 590698 566054
rect 590142 565498 590378 565734
rect 590462 565498 590698 565734
rect 590142 531818 590378 532054
rect 590462 531818 590698 532054
rect 590142 531498 590378 531734
rect 590462 531498 590698 531734
rect 590142 497818 590378 498054
rect 590462 497818 590698 498054
rect 590142 497498 590378 497734
rect 590462 497498 590698 497734
rect 590142 463818 590378 464054
rect 590462 463818 590698 464054
rect 590142 463498 590378 463734
rect 590462 463498 590698 463734
rect 590142 429818 590378 430054
rect 590462 429818 590698 430054
rect 590142 429498 590378 429734
rect 590462 429498 590698 429734
rect 590142 395818 590378 396054
rect 590462 395818 590698 396054
rect 590142 395498 590378 395734
rect 590462 395498 590698 395734
rect 590142 361818 590378 362054
rect 590462 361818 590698 362054
rect 590142 361498 590378 361734
rect 590462 361498 590698 361734
rect 590142 327818 590378 328054
rect 590462 327818 590698 328054
rect 590142 327498 590378 327734
rect 590462 327498 590698 327734
rect 590142 293818 590378 294054
rect 590462 293818 590698 294054
rect 590142 293498 590378 293734
rect 590462 293498 590698 293734
rect 590142 259818 590378 260054
rect 590462 259818 590698 260054
rect 590142 259498 590378 259734
rect 590462 259498 590698 259734
rect 590142 225818 590378 226054
rect 590462 225818 590698 226054
rect 590142 225498 590378 225734
rect 590462 225498 590698 225734
rect 590142 191818 590378 192054
rect 590462 191818 590698 192054
rect 590142 191498 590378 191734
rect 590462 191498 590698 191734
rect 590142 157818 590378 158054
rect 590462 157818 590698 158054
rect 590142 157498 590378 157734
rect 590462 157498 590698 157734
rect 590142 123818 590378 124054
rect 590462 123818 590698 124054
rect 590142 123498 590378 123734
rect 590462 123498 590698 123734
rect 590142 89818 590378 90054
rect 590462 89818 590698 90054
rect 590142 89498 590378 89734
rect 590462 89498 590698 89734
rect 590142 55818 590378 56054
rect 590462 55818 590698 56054
rect 590142 55498 590378 55734
rect 590462 55498 590698 55734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 671538 591338 671774
rect 591422 671538 591658 671774
rect 591102 671218 591338 671454
rect 591422 671218 591658 671454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 603538 591338 603774
rect 591422 603538 591658 603774
rect 591102 603218 591338 603454
rect 591422 603218 591658 603454
rect 591102 569538 591338 569774
rect 591422 569538 591658 569774
rect 591102 569218 591338 569454
rect 591422 569218 591658 569454
rect 591102 535538 591338 535774
rect 591422 535538 591658 535774
rect 591102 535218 591338 535454
rect 591422 535218 591658 535454
rect 591102 501538 591338 501774
rect 591422 501538 591658 501774
rect 591102 501218 591338 501454
rect 591422 501218 591658 501454
rect 591102 467538 591338 467774
rect 591422 467538 591658 467774
rect 591102 467218 591338 467454
rect 591422 467218 591658 467454
rect 591102 433538 591338 433774
rect 591422 433538 591658 433774
rect 591102 433218 591338 433454
rect 591422 433218 591658 433454
rect 591102 399538 591338 399774
rect 591422 399538 591658 399774
rect 591102 399218 591338 399454
rect 591422 399218 591658 399454
rect 591102 365538 591338 365774
rect 591422 365538 591658 365774
rect 591102 365218 591338 365454
rect 591422 365218 591658 365454
rect 591102 331538 591338 331774
rect 591422 331538 591658 331774
rect 591102 331218 591338 331454
rect 591422 331218 591658 331454
rect 591102 297538 591338 297774
rect 591422 297538 591658 297774
rect 591102 297218 591338 297454
rect 591422 297218 591658 297454
rect 591102 263538 591338 263774
rect 591422 263538 591658 263774
rect 591102 263218 591338 263454
rect 591422 263218 591658 263454
rect 591102 229538 591338 229774
rect 591422 229538 591658 229774
rect 591102 229218 591338 229454
rect 591422 229218 591658 229454
rect 591102 195538 591338 195774
rect 591422 195538 591658 195774
rect 591102 195218 591338 195454
rect 591422 195218 591658 195454
rect 591102 161538 591338 161774
rect 591422 161538 591658 161774
rect 591102 161218 591338 161454
rect 591422 161218 591658 161454
rect 591102 127538 591338 127774
rect 591422 127538 591658 127774
rect 591102 127218 591338 127454
rect 591422 127218 591658 127454
rect 591102 93538 591338 93774
rect 591422 93538 591658 93774
rect 591102 93218 591338 93454
rect 591422 93218 591658 93454
rect 591102 59538 591338 59774
rect 591422 59538 591658 59774
rect 591102 59218 591338 59454
rect 591422 59218 591658 59454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 675258 592298 675494
rect 592382 675258 592618 675494
rect 592062 674938 592298 675174
rect 592382 674938 592618 675174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 607258 592298 607494
rect 592382 607258 592618 607494
rect 592062 606938 592298 607174
rect 592382 606938 592618 607174
rect 592062 573258 592298 573494
rect 592382 573258 592618 573494
rect 592062 572938 592298 573174
rect 592382 572938 592618 573174
rect 592062 539258 592298 539494
rect 592382 539258 592618 539494
rect 592062 538938 592298 539174
rect 592382 538938 592618 539174
rect 592062 505258 592298 505494
rect 592382 505258 592618 505494
rect 592062 504938 592298 505174
rect 592382 504938 592618 505174
rect 592062 471258 592298 471494
rect 592382 471258 592618 471494
rect 592062 470938 592298 471174
rect 592382 470938 592618 471174
rect 592062 437258 592298 437494
rect 592382 437258 592618 437494
rect 592062 436938 592298 437174
rect 592382 436938 592618 437174
rect 592062 403258 592298 403494
rect 592382 403258 592618 403494
rect 592062 402938 592298 403174
rect 592382 402938 592618 403174
rect 592062 369258 592298 369494
rect 592382 369258 592618 369494
rect 592062 368938 592298 369174
rect 592382 368938 592618 369174
rect 592062 335258 592298 335494
rect 592382 335258 592618 335494
rect 592062 334938 592298 335174
rect 592382 334938 592618 335174
rect 592062 301258 592298 301494
rect 592382 301258 592618 301494
rect 592062 300938 592298 301174
rect 592382 300938 592618 301174
rect 592062 267258 592298 267494
rect 592382 267258 592618 267494
rect 592062 266938 592298 267174
rect 592382 266938 592618 267174
rect 592062 233258 592298 233494
rect 592382 233258 592618 233494
rect 592062 232938 592298 233174
rect 592382 232938 592618 233174
rect 592062 199258 592298 199494
rect 592382 199258 592618 199494
rect 592062 198938 592298 199174
rect 592382 198938 592618 199174
rect 592062 165258 592298 165494
rect 592382 165258 592618 165494
rect 592062 164938 592298 165174
rect 592382 164938 592618 165174
rect 592062 131258 592298 131494
rect 592382 131258 592618 131494
rect 592062 130938 592298 131174
rect 592382 130938 592618 131174
rect 592062 97258 592298 97494
rect 592382 97258 592618 97494
rect 592062 96938 592298 97174
rect 592382 96938 592618 97174
rect 592062 63258 592298 63494
rect 592382 63258 592618 63494
rect 592062 62938 592298 63174
rect 592382 62938 592618 63174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 61866 711558
rect 62102 711322 62186 711558
rect 62422 711322 95866 711558
rect 96102 711322 96186 711558
rect 96422 711322 129866 711558
rect 130102 711322 130186 711558
rect 130422 711322 163866 711558
rect 164102 711322 164186 711558
rect 164422 711322 197866 711558
rect 198102 711322 198186 711558
rect 198422 711322 231866 711558
rect 232102 711322 232186 711558
rect 232422 711322 265866 711558
rect 266102 711322 266186 711558
rect 266422 711322 299866 711558
rect 300102 711322 300186 711558
rect 300422 711322 333866 711558
rect 334102 711322 334186 711558
rect 334422 711322 367866 711558
rect 368102 711322 368186 711558
rect 368422 711322 401866 711558
rect 402102 711322 402186 711558
rect 402422 711322 435866 711558
rect 436102 711322 436186 711558
rect 436422 711322 469866 711558
rect 470102 711322 470186 711558
rect 470422 711322 503866 711558
rect 504102 711322 504186 711558
rect 504422 711322 537866 711558
rect 538102 711322 538186 711558
rect 538422 711322 571866 711558
rect 572102 711322 572186 711558
rect 572422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 61866 711238
rect 62102 711002 62186 711238
rect 62422 711002 95866 711238
rect 96102 711002 96186 711238
rect 96422 711002 129866 711238
rect 130102 711002 130186 711238
rect 130422 711002 163866 711238
rect 164102 711002 164186 711238
rect 164422 711002 197866 711238
rect 198102 711002 198186 711238
rect 198422 711002 231866 711238
rect 232102 711002 232186 711238
rect 232422 711002 265866 711238
rect 266102 711002 266186 711238
rect 266422 711002 299866 711238
rect 300102 711002 300186 711238
rect 300422 711002 333866 711238
rect 334102 711002 334186 711238
rect 334422 711002 367866 711238
rect 368102 711002 368186 711238
rect 368422 711002 401866 711238
rect 402102 711002 402186 711238
rect 402422 711002 435866 711238
rect 436102 711002 436186 711238
rect 436422 711002 469866 711238
rect 470102 711002 470186 711238
rect 470422 711002 503866 711238
rect 504102 711002 504186 711238
rect 504422 711002 537866 711238
rect 538102 711002 538186 711238
rect 538422 711002 571866 711238
rect 572102 711002 572186 711238
rect 572422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 58146 710598
rect 58382 710362 58466 710598
rect 58702 710362 92146 710598
rect 92382 710362 92466 710598
rect 92702 710362 126146 710598
rect 126382 710362 126466 710598
rect 126702 710362 160146 710598
rect 160382 710362 160466 710598
rect 160702 710362 194146 710598
rect 194382 710362 194466 710598
rect 194702 710362 228146 710598
rect 228382 710362 228466 710598
rect 228702 710362 262146 710598
rect 262382 710362 262466 710598
rect 262702 710362 296146 710598
rect 296382 710362 296466 710598
rect 296702 710362 330146 710598
rect 330382 710362 330466 710598
rect 330702 710362 364146 710598
rect 364382 710362 364466 710598
rect 364702 710362 398146 710598
rect 398382 710362 398466 710598
rect 398702 710362 432146 710598
rect 432382 710362 432466 710598
rect 432702 710362 466146 710598
rect 466382 710362 466466 710598
rect 466702 710362 500146 710598
rect 500382 710362 500466 710598
rect 500702 710362 534146 710598
rect 534382 710362 534466 710598
rect 534702 710362 568146 710598
rect 568382 710362 568466 710598
rect 568702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 58146 710278
rect 58382 710042 58466 710278
rect 58702 710042 92146 710278
rect 92382 710042 92466 710278
rect 92702 710042 126146 710278
rect 126382 710042 126466 710278
rect 126702 710042 160146 710278
rect 160382 710042 160466 710278
rect 160702 710042 194146 710278
rect 194382 710042 194466 710278
rect 194702 710042 228146 710278
rect 228382 710042 228466 710278
rect 228702 710042 262146 710278
rect 262382 710042 262466 710278
rect 262702 710042 296146 710278
rect 296382 710042 296466 710278
rect 296702 710042 330146 710278
rect 330382 710042 330466 710278
rect 330702 710042 364146 710278
rect 364382 710042 364466 710278
rect 364702 710042 398146 710278
rect 398382 710042 398466 710278
rect 398702 710042 432146 710278
rect 432382 710042 432466 710278
rect 432702 710042 466146 710278
rect 466382 710042 466466 710278
rect 466702 710042 500146 710278
rect 500382 710042 500466 710278
rect 500702 710042 534146 710278
rect 534382 710042 534466 710278
rect 534702 710042 568146 710278
rect 568382 710042 568466 710278
rect 568702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 54426 709638
rect 54662 709402 54746 709638
rect 54982 709402 88426 709638
rect 88662 709402 88746 709638
rect 88982 709402 122426 709638
rect 122662 709402 122746 709638
rect 122982 709402 156426 709638
rect 156662 709402 156746 709638
rect 156982 709402 190426 709638
rect 190662 709402 190746 709638
rect 190982 709402 224426 709638
rect 224662 709402 224746 709638
rect 224982 709402 258426 709638
rect 258662 709402 258746 709638
rect 258982 709402 292426 709638
rect 292662 709402 292746 709638
rect 292982 709402 326426 709638
rect 326662 709402 326746 709638
rect 326982 709402 360426 709638
rect 360662 709402 360746 709638
rect 360982 709402 394426 709638
rect 394662 709402 394746 709638
rect 394982 709402 428426 709638
rect 428662 709402 428746 709638
rect 428982 709402 462426 709638
rect 462662 709402 462746 709638
rect 462982 709402 496426 709638
rect 496662 709402 496746 709638
rect 496982 709402 530426 709638
rect 530662 709402 530746 709638
rect 530982 709402 564426 709638
rect 564662 709402 564746 709638
rect 564982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 54426 709318
rect 54662 709082 54746 709318
rect 54982 709082 88426 709318
rect 88662 709082 88746 709318
rect 88982 709082 122426 709318
rect 122662 709082 122746 709318
rect 122982 709082 156426 709318
rect 156662 709082 156746 709318
rect 156982 709082 190426 709318
rect 190662 709082 190746 709318
rect 190982 709082 224426 709318
rect 224662 709082 224746 709318
rect 224982 709082 258426 709318
rect 258662 709082 258746 709318
rect 258982 709082 292426 709318
rect 292662 709082 292746 709318
rect 292982 709082 326426 709318
rect 326662 709082 326746 709318
rect 326982 709082 360426 709318
rect 360662 709082 360746 709318
rect 360982 709082 394426 709318
rect 394662 709082 394746 709318
rect 394982 709082 428426 709318
rect 428662 709082 428746 709318
rect 428982 709082 462426 709318
rect 462662 709082 462746 709318
rect 462982 709082 496426 709318
rect 496662 709082 496746 709318
rect 496982 709082 530426 709318
rect 530662 709082 530746 709318
rect 530982 709082 564426 709318
rect 564662 709082 564746 709318
rect 564982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 50706 708678
rect 50942 708442 51026 708678
rect 51262 708442 84706 708678
rect 84942 708442 85026 708678
rect 85262 708442 118706 708678
rect 118942 708442 119026 708678
rect 119262 708442 152706 708678
rect 152942 708442 153026 708678
rect 153262 708442 186706 708678
rect 186942 708442 187026 708678
rect 187262 708442 220706 708678
rect 220942 708442 221026 708678
rect 221262 708442 254706 708678
rect 254942 708442 255026 708678
rect 255262 708442 288706 708678
rect 288942 708442 289026 708678
rect 289262 708442 322706 708678
rect 322942 708442 323026 708678
rect 323262 708442 356706 708678
rect 356942 708442 357026 708678
rect 357262 708442 390706 708678
rect 390942 708442 391026 708678
rect 391262 708442 424706 708678
rect 424942 708442 425026 708678
rect 425262 708442 458706 708678
rect 458942 708442 459026 708678
rect 459262 708442 492706 708678
rect 492942 708442 493026 708678
rect 493262 708442 526706 708678
rect 526942 708442 527026 708678
rect 527262 708442 560706 708678
rect 560942 708442 561026 708678
rect 561262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 50706 708358
rect 50942 708122 51026 708358
rect 51262 708122 84706 708358
rect 84942 708122 85026 708358
rect 85262 708122 118706 708358
rect 118942 708122 119026 708358
rect 119262 708122 152706 708358
rect 152942 708122 153026 708358
rect 153262 708122 186706 708358
rect 186942 708122 187026 708358
rect 187262 708122 220706 708358
rect 220942 708122 221026 708358
rect 221262 708122 254706 708358
rect 254942 708122 255026 708358
rect 255262 708122 288706 708358
rect 288942 708122 289026 708358
rect 289262 708122 322706 708358
rect 322942 708122 323026 708358
rect 323262 708122 356706 708358
rect 356942 708122 357026 708358
rect 357262 708122 390706 708358
rect 390942 708122 391026 708358
rect 391262 708122 424706 708358
rect 424942 708122 425026 708358
rect 425262 708122 458706 708358
rect 458942 708122 459026 708358
rect 459262 708122 492706 708358
rect 492942 708122 493026 708358
rect 493262 708122 526706 708358
rect 526942 708122 527026 708358
rect 527262 708122 560706 708358
rect 560942 708122 561026 708358
rect 561262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 46986 707718
rect 47222 707482 47306 707718
rect 47542 707482 80986 707718
rect 81222 707482 81306 707718
rect 81542 707482 114986 707718
rect 115222 707482 115306 707718
rect 115542 707482 148986 707718
rect 149222 707482 149306 707718
rect 149542 707482 182986 707718
rect 183222 707482 183306 707718
rect 183542 707482 216986 707718
rect 217222 707482 217306 707718
rect 217542 707482 250986 707718
rect 251222 707482 251306 707718
rect 251542 707482 284986 707718
rect 285222 707482 285306 707718
rect 285542 707482 318986 707718
rect 319222 707482 319306 707718
rect 319542 707482 352986 707718
rect 353222 707482 353306 707718
rect 353542 707482 386986 707718
rect 387222 707482 387306 707718
rect 387542 707482 420986 707718
rect 421222 707482 421306 707718
rect 421542 707482 454986 707718
rect 455222 707482 455306 707718
rect 455542 707482 488986 707718
rect 489222 707482 489306 707718
rect 489542 707482 522986 707718
rect 523222 707482 523306 707718
rect 523542 707482 556986 707718
rect 557222 707482 557306 707718
rect 557542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 46986 707398
rect 47222 707162 47306 707398
rect 47542 707162 80986 707398
rect 81222 707162 81306 707398
rect 81542 707162 114986 707398
rect 115222 707162 115306 707398
rect 115542 707162 148986 707398
rect 149222 707162 149306 707398
rect 149542 707162 182986 707398
rect 183222 707162 183306 707398
rect 183542 707162 216986 707398
rect 217222 707162 217306 707398
rect 217542 707162 250986 707398
rect 251222 707162 251306 707398
rect 251542 707162 284986 707398
rect 285222 707162 285306 707398
rect 285542 707162 318986 707398
rect 319222 707162 319306 707398
rect 319542 707162 352986 707398
rect 353222 707162 353306 707398
rect 353542 707162 386986 707398
rect 387222 707162 387306 707398
rect 387542 707162 420986 707398
rect 421222 707162 421306 707398
rect 421542 707162 454986 707398
rect 455222 707162 455306 707398
rect 455542 707162 488986 707398
rect 489222 707162 489306 707398
rect 489542 707162 522986 707398
rect 523222 707162 523306 707398
rect 523542 707162 556986 707398
rect 557222 707162 557306 707398
rect 557542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 43266 706758
rect 43502 706522 43586 706758
rect 43822 706522 77266 706758
rect 77502 706522 77586 706758
rect 77822 706522 111266 706758
rect 111502 706522 111586 706758
rect 111822 706522 145266 706758
rect 145502 706522 145586 706758
rect 145822 706522 179266 706758
rect 179502 706522 179586 706758
rect 179822 706522 213266 706758
rect 213502 706522 213586 706758
rect 213822 706522 247266 706758
rect 247502 706522 247586 706758
rect 247822 706522 281266 706758
rect 281502 706522 281586 706758
rect 281822 706522 315266 706758
rect 315502 706522 315586 706758
rect 315822 706522 349266 706758
rect 349502 706522 349586 706758
rect 349822 706522 383266 706758
rect 383502 706522 383586 706758
rect 383822 706522 417266 706758
rect 417502 706522 417586 706758
rect 417822 706522 451266 706758
rect 451502 706522 451586 706758
rect 451822 706522 485266 706758
rect 485502 706522 485586 706758
rect 485822 706522 519266 706758
rect 519502 706522 519586 706758
rect 519822 706522 553266 706758
rect 553502 706522 553586 706758
rect 553822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 43266 706438
rect 43502 706202 43586 706438
rect 43822 706202 77266 706438
rect 77502 706202 77586 706438
rect 77822 706202 111266 706438
rect 111502 706202 111586 706438
rect 111822 706202 145266 706438
rect 145502 706202 145586 706438
rect 145822 706202 179266 706438
rect 179502 706202 179586 706438
rect 179822 706202 213266 706438
rect 213502 706202 213586 706438
rect 213822 706202 247266 706438
rect 247502 706202 247586 706438
rect 247822 706202 281266 706438
rect 281502 706202 281586 706438
rect 281822 706202 315266 706438
rect 315502 706202 315586 706438
rect 315822 706202 349266 706438
rect 349502 706202 349586 706438
rect 349822 706202 383266 706438
rect 383502 706202 383586 706438
rect 383822 706202 417266 706438
rect 417502 706202 417586 706438
rect 417822 706202 451266 706438
rect 451502 706202 451586 706438
rect 451822 706202 485266 706438
rect 485502 706202 485586 706438
rect 485822 706202 519266 706438
rect 519502 706202 519586 706438
rect 519822 706202 553266 706438
rect 553502 706202 553586 706438
rect 553822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 39546 705798
rect 39782 705562 39866 705798
rect 40102 705562 73546 705798
rect 73782 705562 73866 705798
rect 74102 705562 107546 705798
rect 107782 705562 107866 705798
rect 108102 705562 141546 705798
rect 141782 705562 141866 705798
rect 142102 705562 175546 705798
rect 175782 705562 175866 705798
rect 176102 705562 209546 705798
rect 209782 705562 209866 705798
rect 210102 705562 243546 705798
rect 243782 705562 243866 705798
rect 244102 705562 277546 705798
rect 277782 705562 277866 705798
rect 278102 705562 311546 705798
rect 311782 705562 311866 705798
rect 312102 705562 345546 705798
rect 345782 705562 345866 705798
rect 346102 705562 379546 705798
rect 379782 705562 379866 705798
rect 380102 705562 413546 705798
rect 413782 705562 413866 705798
rect 414102 705562 447546 705798
rect 447782 705562 447866 705798
rect 448102 705562 481546 705798
rect 481782 705562 481866 705798
rect 482102 705562 515546 705798
rect 515782 705562 515866 705798
rect 516102 705562 549546 705798
rect 549782 705562 549866 705798
rect 550102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 39546 705478
rect 39782 705242 39866 705478
rect 40102 705242 73546 705478
rect 73782 705242 73866 705478
rect 74102 705242 107546 705478
rect 107782 705242 107866 705478
rect 108102 705242 141546 705478
rect 141782 705242 141866 705478
rect 142102 705242 175546 705478
rect 175782 705242 175866 705478
rect 176102 705242 209546 705478
rect 209782 705242 209866 705478
rect 210102 705242 243546 705478
rect 243782 705242 243866 705478
rect 244102 705242 277546 705478
rect 277782 705242 277866 705478
rect 278102 705242 311546 705478
rect 311782 705242 311866 705478
rect 312102 705242 345546 705478
rect 345782 705242 345866 705478
rect 346102 705242 379546 705478
rect 379782 705242 379866 705478
rect 380102 705242 413546 705478
rect 413782 705242 413866 705478
rect 414102 705242 447546 705478
rect 447782 705242 447866 705478
rect 448102 705242 481546 705478
rect 481782 705242 481866 705478
rect 482102 705242 515546 705478
rect 515782 705242 515866 705478
rect 516102 705242 549546 705478
rect 549782 705242 549866 705478
rect 550102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 35826 704838
rect 36062 704602 36146 704838
rect 36382 704602 69826 704838
rect 70062 704602 70146 704838
rect 70382 704602 103826 704838
rect 104062 704602 104146 704838
rect 104382 704602 137826 704838
rect 138062 704602 138146 704838
rect 138382 704602 171826 704838
rect 172062 704602 172146 704838
rect 172382 704602 205826 704838
rect 206062 704602 206146 704838
rect 206382 704602 239826 704838
rect 240062 704602 240146 704838
rect 240382 704602 273826 704838
rect 274062 704602 274146 704838
rect 274382 704602 307826 704838
rect 308062 704602 308146 704838
rect 308382 704602 341826 704838
rect 342062 704602 342146 704838
rect 342382 704602 375826 704838
rect 376062 704602 376146 704838
rect 376382 704602 409826 704838
rect 410062 704602 410146 704838
rect 410382 704602 443826 704838
rect 444062 704602 444146 704838
rect 444382 704602 477826 704838
rect 478062 704602 478146 704838
rect 478382 704602 511826 704838
rect 512062 704602 512146 704838
rect 512382 704602 545826 704838
rect 546062 704602 546146 704838
rect 546382 704602 579826 704838
rect 580062 704602 580146 704838
rect 580382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 35826 704518
rect 36062 704282 36146 704518
rect 36382 704282 69826 704518
rect 70062 704282 70146 704518
rect 70382 704282 103826 704518
rect 104062 704282 104146 704518
rect 104382 704282 137826 704518
rect 138062 704282 138146 704518
rect 138382 704282 171826 704518
rect 172062 704282 172146 704518
rect 172382 704282 205826 704518
rect 206062 704282 206146 704518
rect 206382 704282 239826 704518
rect 240062 704282 240146 704518
rect 240382 704282 273826 704518
rect 274062 704282 274146 704518
rect 274382 704282 307826 704518
rect 308062 704282 308146 704518
rect 308382 704282 341826 704518
rect 342062 704282 342146 704518
rect 342382 704282 375826 704518
rect 376062 704282 376146 704518
rect 376382 704282 409826 704518
rect 410062 704282 410146 704518
rect 410382 704282 443826 704518
rect 444062 704282 444146 704518
rect 444382 704282 477826 704518
rect 478062 704282 478146 704518
rect 478382 704282 511826 704518
rect 512062 704282 512146 704518
rect 512382 704282 545826 704518
rect 546062 704282 546146 704518
rect 546382 704282 579826 704518
rect 580062 704282 580146 704518
rect 580382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698334 592650 698366
rect -8726 698098 -5814 698334
rect -5578 698098 -5494 698334
rect -5258 698098 16706 698334
rect 16942 698098 17026 698334
rect 17262 698098 50706 698334
rect 50942 698098 51026 698334
rect 51262 698098 84706 698334
rect 84942 698098 85026 698334
rect 85262 698098 118706 698334
rect 118942 698098 119026 698334
rect 119262 698098 152706 698334
rect 152942 698098 153026 698334
rect 153262 698098 186706 698334
rect 186942 698098 187026 698334
rect 187262 698098 220706 698334
rect 220942 698098 221026 698334
rect 221262 698098 254706 698334
rect 254942 698098 255026 698334
rect 255262 698098 288706 698334
rect 288942 698098 289026 698334
rect 289262 698098 322706 698334
rect 322942 698098 323026 698334
rect 323262 698098 356706 698334
rect 356942 698098 357026 698334
rect 357262 698098 390706 698334
rect 390942 698098 391026 698334
rect 391262 698098 424706 698334
rect 424942 698098 425026 698334
rect 425262 698098 458706 698334
rect 458942 698098 459026 698334
rect 459262 698098 492706 698334
rect 492942 698098 493026 698334
rect 493262 698098 526706 698334
rect 526942 698098 527026 698334
rect 527262 698098 560706 698334
rect 560942 698098 561026 698334
rect 561262 698098 589182 698334
rect 589418 698098 589502 698334
rect 589738 698098 592650 698334
rect -8726 698014 592650 698098
rect -8726 697778 -5814 698014
rect -5578 697778 -5494 698014
rect -5258 697778 16706 698014
rect 16942 697778 17026 698014
rect 17262 697778 50706 698014
rect 50942 697778 51026 698014
rect 51262 697778 84706 698014
rect 84942 697778 85026 698014
rect 85262 697778 118706 698014
rect 118942 697778 119026 698014
rect 119262 697778 152706 698014
rect 152942 697778 153026 698014
rect 153262 697778 186706 698014
rect 186942 697778 187026 698014
rect 187262 697778 220706 698014
rect 220942 697778 221026 698014
rect 221262 697778 254706 698014
rect 254942 697778 255026 698014
rect 255262 697778 288706 698014
rect 288942 697778 289026 698014
rect 289262 697778 322706 698014
rect 322942 697778 323026 698014
rect 323262 697778 356706 698014
rect 356942 697778 357026 698014
rect 357262 697778 390706 698014
rect 390942 697778 391026 698014
rect 391262 697778 424706 698014
rect 424942 697778 425026 698014
rect 425262 697778 458706 698014
rect 458942 697778 459026 698014
rect 459262 697778 492706 698014
rect 492942 697778 493026 698014
rect 493262 697778 526706 698014
rect 526942 697778 527026 698014
rect 527262 697778 560706 698014
rect 560942 697778 561026 698014
rect 561262 697778 589182 698014
rect 589418 697778 589502 698014
rect 589738 697778 592650 698014
rect -8726 697746 592650 697778
rect -8726 694614 592650 694646
rect -8726 694378 -4854 694614
rect -4618 694378 -4534 694614
rect -4298 694378 12986 694614
rect 13222 694378 13306 694614
rect 13542 694378 46986 694614
rect 47222 694378 47306 694614
rect 47542 694378 80986 694614
rect 81222 694378 81306 694614
rect 81542 694378 114986 694614
rect 115222 694378 115306 694614
rect 115542 694378 148986 694614
rect 149222 694378 149306 694614
rect 149542 694378 182986 694614
rect 183222 694378 183306 694614
rect 183542 694378 216986 694614
rect 217222 694378 217306 694614
rect 217542 694378 250986 694614
rect 251222 694378 251306 694614
rect 251542 694378 284986 694614
rect 285222 694378 285306 694614
rect 285542 694378 318986 694614
rect 319222 694378 319306 694614
rect 319542 694378 352986 694614
rect 353222 694378 353306 694614
rect 353542 694378 386986 694614
rect 387222 694378 387306 694614
rect 387542 694378 420986 694614
rect 421222 694378 421306 694614
rect 421542 694378 454986 694614
rect 455222 694378 455306 694614
rect 455542 694378 488986 694614
rect 489222 694378 489306 694614
rect 489542 694378 522986 694614
rect 523222 694378 523306 694614
rect 523542 694378 556986 694614
rect 557222 694378 557306 694614
rect 557542 694378 588222 694614
rect 588458 694378 588542 694614
rect 588778 694378 592650 694614
rect -8726 694294 592650 694378
rect -8726 694058 -4854 694294
rect -4618 694058 -4534 694294
rect -4298 694058 12986 694294
rect 13222 694058 13306 694294
rect 13542 694058 46986 694294
rect 47222 694058 47306 694294
rect 47542 694058 80986 694294
rect 81222 694058 81306 694294
rect 81542 694058 114986 694294
rect 115222 694058 115306 694294
rect 115542 694058 148986 694294
rect 149222 694058 149306 694294
rect 149542 694058 182986 694294
rect 183222 694058 183306 694294
rect 183542 694058 216986 694294
rect 217222 694058 217306 694294
rect 217542 694058 250986 694294
rect 251222 694058 251306 694294
rect 251542 694058 284986 694294
rect 285222 694058 285306 694294
rect 285542 694058 318986 694294
rect 319222 694058 319306 694294
rect 319542 694058 352986 694294
rect 353222 694058 353306 694294
rect 353542 694058 386986 694294
rect 387222 694058 387306 694294
rect 387542 694058 420986 694294
rect 421222 694058 421306 694294
rect 421542 694058 454986 694294
rect 455222 694058 455306 694294
rect 455542 694058 488986 694294
rect 489222 694058 489306 694294
rect 489542 694058 522986 694294
rect 523222 694058 523306 694294
rect 523542 694058 556986 694294
rect 557222 694058 557306 694294
rect 557542 694058 588222 694294
rect 588458 694058 588542 694294
rect 588778 694058 592650 694294
rect -8726 694026 592650 694058
rect -8726 690894 592650 690926
rect -8726 690658 -3894 690894
rect -3658 690658 -3574 690894
rect -3338 690658 9266 690894
rect 9502 690658 9586 690894
rect 9822 690658 43266 690894
rect 43502 690658 43586 690894
rect 43822 690658 77266 690894
rect 77502 690658 77586 690894
rect 77822 690658 111266 690894
rect 111502 690658 111586 690894
rect 111822 690658 145266 690894
rect 145502 690658 145586 690894
rect 145822 690658 179266 690894
rect 179502 690658 179586 690894
rect 179822 690658 213266 690894
rect 213502 690658 213586 690894
rect 213822 690658 247266 690894
rect 247502 690658 247586 690894
rect 247822 690658 281266 690894
rect 281502 690658 281586 690894
rect 281822 690658 315266 690894
rect 315502 690658 315586 690894
rect 315822 690658 349266 690894
rect 349502 690658 349586 690894
rect 349822 690658 383266 690894
rect 383502 690658 383586 690894
rect 383822 690658 417266 690894
rect 417502 690658 417586 690894
rect 417822 690658 451266 690894
rect 451502 690658 451586 690894
rect 451822 690658 485266 690894
rect 485502 690658 485586 690894
rect 485822 690658 519266 690894
rect 519502 690658 519586 690894
rect 519822 690658 553266 690894
rect 553502 690658 553586 690894
rect 553822 690658 587262 690894
rect 587498 690658 587582 690894
rect 587818 690658 592650 690894
rect -8726 690574 592650 690658
rect -8726 690338 -3894 690574
rect -3658 690338 -3574 690574
rect -3338 690338 9266 690574
rect 9502 690338 9586 690574
rect 9822 690338 43266 690574
rect 43502 690338 43586 690574
rect 43822 690338 77266 690574
rect 77502 690338 77586 690574
rect 77822 690338 111266 690574
rect 111502 690338 111586 690574
rect 111822 690338 145266 690574
rect 145502 690338 145586 690574
rect 145822 690338 179266 690574
rect 179502 690338 179586 690574
rect 179822 690338 213266 690574
rect 213502 690338 213586 690574
rect 213822 690338 247266 690574
rect 247502 690338 247586 690574
rect 247822 690338 281266 690574
rect 281502 690338 281586 690574
rect 281822 690338 315266 690574
rect 315502 690338 315586 690574
rect 315822 690338 349266 690574
rect 349502 690338 349586 690574
rect 349822 690338 383266 690574
rect 383502 690338 383586 690574
rect 383822 690338 417266 690574
rect 417502 690338 417586 690574
rect 417822 690338 451266 690574
rect 451502 690338 451586 690574
rect 451822 690338 485266 690574
rect 485502 690338 485586 690574
rect 485822 690338 519266 690574
rect 519502 690338 519586 690574
rect 519822 690338 553266 690574
rect 553502 690338 553586 690574
rect 553822 690338 587262 690574
rect 587498 690338 587582 690574
rect 587818 690338 592650 690574
rect -8726 690306 592650 690338
rect -8726 687174 592650 687206
rect -8726 686938 -2934 687174
rect -2698 686938 -2614 687174
rect -2378 686938 5546 687174
rect 5782 686938 5866 687174
rect 6102 686938 39546 687174
rect 39782 686938 39866 687174
rect 40102 686938 73546 687174
rect 73782 686938 73866 687174
rect 74102 686938 107546 687174
rect 107782 686938 107866 687174
rect 108102 686938 141546 687174
rect 141782 686938 141866 687174
rect 142102 686938 175546 687174
rect 175782 686938 175866 687174
rect 176102 686938 209546 687174
rect 209782 686938 209866 687174
rect 210102 686938 243546 687174
rect 243782 686938 243866 687174
rect 244102 686938 277546 687174
rect 277782 686938 277866 687174
rect 278102 686938 311546 687174
rect 311782 686938 311866 687174
rect 312102 686938 345546 687174
rect 345782 686938 345866 687174
rect 346102 686938 379546 687174
rect 379782 686938 379866 687174
rect 380102 686938 413546 687174
rect 413782 686938 413866 687174
rect 414102 686938 447546 687174
rect 447782 686938 447866 687174
rect 448102 686938 481546 687174
rect 481782 686938 481866 687174
rect 482102 686938 515546 687174
rect 515782 686938 515866 687174
rect 516102 686938 549546 687174
rect 549782 686938 549866 687174
rect 550102 686938 586302 687174
rect 586538 686938 586622 687174
rect 586858 686938 592650 687174
rect -8726 686854 592650 686938
rect -8726 686618 -2934 686854
rect -2698 686618 -2614 686854
rect -2378 686618 5546 686854
rect 5782 686618 5866 686854
rect 6102 686618 39546 686854
rect 39782 686618 39866 686854
rect 40102 686618 73546 686854
rect 73782 686618 73866 686854
rect 74102 686618 107546 686854
rect 107782 686618 107866 686854
rect 108102 686618 141546 686854
rect 141782 686618 141866 686854
rect 142102 686618 175546 686854
rect 175782 686618 175866 686854
rect 176102 686618 209546 686854
rect 209782 686618 209866 686854
rect 210102 686618 243546 686854
rect 243782 686618 243866 686854
rect 244102 686618 277546 686854
rect 277782 686618 277866 686854
rect 278102 686618 311546 686854
rect 311782 686618 311866 686854
rect 312102 686618 345546 686854
rect 345782 686618 345866 686854
rect 346102 686618 379546 686854
rect 379782 686618 379866 686854
rect 380102 686618 413546 686854
rect 413782 686618 413866 686854
rect 414102 686618 447546 686854
rect 447782 686618 447866 686854
rect 448102 686618 481546 686854
rect 481782 686618 481866 686854
rect 482102 686618 515546 686854
rect 515782 686618 515866 686854
rect 516102 686618 549546 686854
rect 549782 686618 549866 686854
rect 550102 686618 586302 686854
rect 586538 686618 586622 686854
rect 586858 686618 592650 686854
rect -8726 686586 592650 686618
rect -8726 683454 592650 683486
rect -8726 683218 -1974 683454
rect -1738 683218 -1654 683454
rect -1418 683218 1826 683454
rect 2062 683218 2146 683454
rect 2382 683218 35826 683454
rect 36062 683218 36146 683454
rect 36382 683218 69826 683454
rect 70062 683218 70146 683454
rect 70382 683218 103826 683454
rect 104062 683218 104146 683454
rect 104382 683218 137826 683454
rect 138062 683218 138146 683454
rect 138382 683218 171826 683454
rect 172062 683218 172146 683454
rect 172382 683218 205826 683454
rect 206062 683218 206146 683454
rect 206382 683218 239826 683454
rect 240062 683218 240146 683454
rect 240382 683218 273826 683454
rect 274062 683218 274146 683454
rect 274382 683218 307826 683454
rect 308062 683218 308146 683454
rect 308382 683218 341826 683454
rect 342062 683218 342146 683454
rect 342382 683218 375826 683454
rect 376062 683218 376146 683454
rect 376382 683218 409826 683454
rect 410062 683218 410146 683454
rect 410382 683218 443826 683454
rect 444062 683218 444146 683454
rect 444382 683218 477826 683454
rect 478062 683218 478146 683454
rect 478382 683218 511826 683454
rect 512062 683218 512146 683454
rect 512382 683218 545826 683454
rect 546062 683218 546146 683454
rect 546382 683218 579826 683454
rect 580062 683218 580146 683454
rect 580382 683218 585342 683454
rect 585578 683218 585662 683454
rect 585898 683218 592650 683454
rect -8726 683134 592650 683218
rect -8726 682898 -1974 683134
rect -1738 682898 -1654 683134
rect -1418 682898 1826 683134
rect 2062 682898 2146 683134
rect 2382 682898 35826 683134
rect 36062 682898 36146 683134
rect 36382 682898 69826 683134
rect 70062 682898 70146 683134
rect 70382 682898 103826 683134
rect 104062 682898 104146 683134
rect 104382 682898 137826 683134
rect 138062 682898 138146 683134
rect 138382 682898 171826 683134
rect 172062 682898 172146 683134
rect 172382 682898 205826 683134
rect 206062 682898 206146 683134
rect 206382 682898 239826 683134
rect 240062 682898 240146 683134
rect 240382 682898 273826 683134
rect 274062 682898 274146 683134
rect 274382 682898 307826 683134
rect 308062 682898 308146 683134
rect 308382 682898 341826 683134
rect 342062 682898 342146 683134
rect 342382 682898 375826 683134
rect 376062 682898 376146 683134
rect 376382 682898 409826 683134
rect 410062 682898 410146 683134
rect 410382 682898 443826 683134
rect 444062 682898 444146 683134
rect 444382 682898 477826 683134
rect 478062 682898 478146 683134
rect 478382 682898 511826 683134
rect 512062 682898 512146 683134
rect 512382 682898 545826 683134
rect 546062 682898 546146 683134
rect 546382 682898 579826 683134
rect 580062 682898 580146 683134
rect 580382 682898 585342 683134
rect 585578 682898 585662 683134
rect 585898 682898 592650 683134
rect -8726 682866 592650 682898
rect -8726 675494 592650 675526
rect -8726 675258 -8694 675494
rect -8458 675258 -8374 675494
rect -8138 675258 27866 675494
rect 28102 675258 28186 675494
rect 28422 675258 61866 675494
rect 62102 675258 62186 675494
rect 62422 675258 95866 675494
rect 96102 675258 96186 675494
rect 96422 675258 129866 675494
rect 130102 675258 130186 675494
rect 130422 675258 163866 675494
rect 164102 675258 164186 675494
rect 164422 675258 197866 675494
rect 198102 675258 198186 675494
rect 198422 675258 231866 675494
rect 232102 675258 232186 675494
rect 232422 675258 265866 675494
rect 266102 675258 266186 675494
rect 266422 675258 299866 675494
rect 300102 675258 300186 675494
rect 300422 675258 333866 675494
rect 334102 675258 334186 675494
rect 334422 675258 367866 675494
rect 368102 675258 368186 675494
rect 368422 675258 401866 675494
rect 402102 675258 402186 675494
rect 402422 675258 435866 675494
rect 436102 675258 436186 675494
rect 436422 675258 469866 675494
rect 470102 675258 470186 675494
rect 470422 675258 503866 675494
rect 504102 675258 504186 675494
rect 504422 675258 537866 675494
rect 538102 675258 538186 675494
rect 538422 675258 571866 675494
rect 572102 675258 572186 675494
rect 572422 675258 592062 675494
rect 592298 675258 592382 675494
rect 592618 675258 592650 675494
rect -8726 675174 592650 675258
rect -8726 674938 -8694 675174
rect -8458 674938 -8374 675174
rect -8138 674938 27866 675174
rect 28102 674938 28186 675174
rect 28422 674938 61866 675174
rect 62102 674938 62186 675174
rect 62422 674938 95866 675174
rect 96102 674938 96186 675174
rect 96422 674938 129866 675174
rect 130102 674938 130186 675174
rect 130422 674938 163866 675174
rect 164102 674938 164186 675174
rect 164422 674938 197866 675174
rect 198102 674938 198186 675174
rect 198422 674938 231866 675174
rect 232102 674938 232186 675174
rect 232422 674938 265866 675174
rect 266102 674938 266186 675174
rect 266422 674938 299866 675174
rect 300102 674938 300186 675174
rect 300422 674938 333866 675174
rect 334102 674938 334186 675174
rect 334422 674938 367866 675174
rect 368102 674938 368186 675174
rect 368422 674938 401866 675174
rect 402102 674938 402186 675174
rect 402422 674938 435866 675174
rect 436102 674938 436186 675174
rect 436422 674938 469866 675174
rect 470102 674938 470186 675174
rect 470422 674938 503866 675174
rect 504102 674938 504186 675174
rect 504422 674938 537866 675174
rect 538102 674938 538186 675174
rect 538422 674938 571866 675174
rect 572102 674938 572186 675174
rect 572422 674938 592062 675174
rect 592298 674938 592382 675174
rect 592618 674938 592650 675174
rect -8726 674906 592650 674938
rect -8726 671774 592650 671806
rect -8726 671538 -7734 671774
rect -7498 671538 -7414 671774
rect -7178 671538 24146 671774
rect 24382 671538 24466 671774
rect 24702 671538 58146 671774
rect 58382 671538 58466 671774
rect 58702 671538 92146 671774
rect 92382 671538 92466 671774
rect 92702 671538 126146 671774
rect 126382 671538 126466 671774
rect 126702 671538 160146 671774
rect 160382 671538 160466 671774
rect 160702 671538 194146 671774
rect 194382 671538 194466 671774
rect 194702 671538 228146 671774
rect 228382 671538 228466 671774
rect 228702 671538 262146 671774
rect 262382 671538 262466 671774
rect 262702 671538 296146 671774
rect 296382 671538 296466 671774
rect 296702 671538 330146 671774
rect 330382 671538 330466 671774
rect 330702 671538 364146 671774
rect 364382 671538 364466 671774
rect 364702 671538 398146 671774
rect 398382 671538 398466 671774
rect 398702 671538 432146 671774
rect 432382 671538 432466 671774
rect 432702 671538 466146 671774
rect 466382 671538 466466 671774
rect 466702 671538 500146 671774
rect 500382 671538 500466 671774
rect 500702 671538 534146 671774
rect 534382 671538 534466 671774
rect 534702 671538 568146 671774
rect 568382 671538 568466 671774
rect 568702 671538 591102 671774
rect 591338 671538 591422 671774
rect 591658 671538 592650 671774
rect -8726 671454 592650 671538
rect -8726 671218 -7734 671454
rect -7498 671218 -7414 671454
rect -7178 671218 24146 671454
rect 24382 671218 24466 671454
rect 24702 671218 58146 671454
rect 58382 671218 58466 671454
rect 58702 671218 92146 671454
rect 92382 671218 92466 671454
rect 92702 671218 126146 671454
rect 126382 671218 126466 671454
rect 126702 671218 160146 671454
rect 160382 671218 160466 671454
rect 160702 671218 194146 671454
rect 194382 671218 194466 671454
rect 194702 671218 228146 671454
rect 228382 671218 228466 671454
rect 228702 671218 262146 671454
rect 262382 671218 262466 671454
rect 262702 671218 296146 671454
rect 296382 671218 296466 671454
rect 296702 671218 330146 671454
rect 330382 671218 330466 671454
rect 330702 671218 364146 671454
rect 364382 671218 364466 671454
rect 364702 671218 398146 671454
rect 398382 671218 398466 671454
rect 398702 671218 432146 671454
rect 432382 671218 432466 671454
rect 432702 671218 466146 671454
rect 466382 671218 466466 671454
rect 466702 671218 500146 671454
rect 500382 671218 500466 671454
rect 500702 671218 534146 671454
rect 534382 671218 534466 671454
rect 534702 671218 568146 671454
rect 568382 671218 568466 671454
rect 568702 671218 591102 671454
rect 591338 671218 591422 671454
rect 591658 671218 592650 671454
rect -8726 671186 592650 671218
rect -8726 668054 592650 668086
rect -8726 667818 -6774 668054
rect -6538 667818 -6454 668054
rect -6218 667818 20426 668054
rect 20662 667818 20746 668054
rect 20982 667818 54426 668054
rect 54662 667818 54746 668054
rect 54982 667818 88426 668054
rect 88662 667818 88746 668054
rect 88982 667818 122426 668054
rect 122662 667818 122746 668054
rect 122982 667818 156426 668054
rect 156662 667818 156746 668054
rect 156982 667818 190426 668054
rect 190662 667818 190746 668054
rect 190982 667818 224426 668054
rect 224662 667818 224746 668054
rect 224982 667818 258426 668054
rect 258662 667818 258746 668054
rect 258982 667818 292426 668054
rect 292662 667818 292746 668054
rect 292982 667818 326426 668054
rect 326662 667818 326746 668054
rect 326982 667818 360426 668054
rect 360662 667818 360746 668054
rect 360982 667818 394426 668054
rect 394662 667818 394746 668054
rect 394982 667818 428426 668054
rect 428662 667818 428746 668054
rect 428982 667818 462426 668054
rect 462662 667818 462746 668054
rect 462982 667818 496426 668054
rect 496662 667818 496746 668054
rect 496982 667818 530426 668054
rect 530662 667818 530746 668054
rect 530982 667818 564426 668054
rect 564662 667818 564746 668054
rect 564982 667818 590142 668054
rect 590378 667818 590462 668054
rect 590698 667818 592650 668054
rect -8726 667734 592650 667818
rect -8726 667498 -6774 667734
rect -6538 667498 -6454 667734
rect -6218 667498 20426 667734
rect 20662 667498 20746 667734
rect 20982 667498 54426 667734
rect 54662 667498 54746 667734
rect 54982 667498 88426 667734
rect 88662 667498 88746 667734
rect 88982 667498 122426 667734
rect 122662 667498 122746 667734
rect 122982 667498 156426 667734
rect 156662 667498 156746 667734
rect 156982 667498 190426 667734
rect 190662 667498 190746 667734
rect 190982 667498 224426 667734
rect 224662 667498 224746 667734
rect 224982 667498 258426 667734
rect 258662 667498 258746 667734
rect 258982 667498 292426 667734
rect 292662 667498 292746 667734
rect 292982 667498 326426 667734
rect 326662 667498 326746 667734
rect 326982 667498 360426 667734
rect 360662 667498 360746 667734
rect 360982 667498 394426 667734
rect 394662 667498 394746 667734
rect 394982 667498 428426 667734
rect 428662 667498 428746 667734
rect 428982 667498 462426 667734
rect 462662 667498 462746 667734
rect 462982 667498 496426 667734
rect 496662 667498 496746 667734
rect 496982 667498 530426 667734
rect 530662 667498 530746 667734
rect 530982 667498 564426 667734
rect 564662 667498 564746 667734
rect 564982 667498 590142 667734
rect 590378 667498 590462 667734
rect 590698 667498 592650 667734
rect -8726 667466 592650 667498
rect -8726 664334 592650 664366
rect -8726 664098 -5814 664334
rect -5578 664098 -5494 664334
rect -5258 664098 16706 664334
rect 16942 664098 17026 664334
rect 17262 664098 50706 664334
rect 50942 664098 51026 664334
rect 51262 664098 84706 664334
rect 84942 664098 85026 664334
rect 85262 664098 118706 664334
rect 118942 664098 119026 664334
rect 119262 664098 152706 664334
rect 152942 664098 153026 664334
rect 153262 664098 186706 664334
rect 186942 664098 187026 664334
rect 187262 664098 220706 664334
rect 220942 664098 221026 664334
rect 221262 664098 254706 664334
rect 254942 664098 255026 664334
rect 255262 664098 288706 664334
rect 288942 664098 289026 664334
rect 289262 664098 322706 664334
rect 322942 664098 323026 664334
rect 323262 664098 356706 664334
rect 356942 664098 357026 664334
rect 357262 664098 390706 664334
rect 390942 664098 391026 664334
rect 391262 664098 424706 664334
rect 424942 664098 425026 664334
rect 425262 664098 458706 664334
rect 458942 664098 459026 664334
rect 459262 664098 492706 664334
rect 492942 664098 493026 664334
rect 493262 664098 526706 664334
rect 526942 664098 527026 664334
rect 527262 664098 560706 664334
rect 560942 664098 561026 664334
rect 561262 664098 589182 664334
rect 589418 664098 589502 664334
rect 589738 664098 592650 664334
rect -8726 664014 592650 664098
rect -8726 663778 -5814 664014
rect -5578 663778 -5494 664014
rect -5258 663778 16706 664014
rect 16942 663778 17026 664014
rect 17262 663778 50706 664014
rect 50942 663778 51026 664014
rect 51262 663778 84706 664014
rect 84942 663778 85026 664014
rect 85262 663778 118706 664014
rect 118942 663778 119026 664014
rect 119262 663778 152706 664014
rect 152942 663778 153026 664014
rect 153262 663778 186706 664014
rect 186942 663778 187026 664014
rect 187262 663778 220706 664014
rect 220942 663778 221026 664014
rect 221262 663778 254706 664014
rect 254942 663778 255026 664014
rect 255262 663778 288706 664014
rect 288942 663778 289026 664014
rect 289262 663778 322706 664014
rect 322942 663778 323026 664014
rect 323262 663778 356706 664014
rect 356942 663778 357026 664014
rect 357262 663778 390706 664014
rect 390942 663778 391026 664014
rect 391262 663778 424706 664014
rect 424942 663778 425026 664014
rect 425262 663778 458706 664014
rect 458942 663778 459026 664014
rect 459262 663778 492706 664014
rect 492942 663778 493026 664014
rect 493262 663778 526706 664014
rect 526942 663778 527026 664014
rect 527262 663778 560706 664014
rect 560942 663778 561026 664014
rect 561262 663778 589182 664014
rect 589418 663778 589502 664014
rect 589738 663778 592650 664014
rect -8726 663746 592650 663778
rect -8726 660614 592650 660646
rect -8726 660378 -4854 660614
rect -4618 660378 -4534 660614
rect -4298 660378 12986 660614
rect 13222 660378 13306 660614
rect 13542 660378 46986 660614
rect 47222 660378 47306 660614
rect 47542 660378 80986 660614
rect 81222 660378 81306 660614
rect 81542 660378 114986 660614
rect 115222 660378 115306 660614
rect 115542 660378 148986 660614
rect 149222 660378 149306 660614
rect 149542 660378 182986 660614
rect 183222 660378 183306 660614
rect 183542 660378 216986 660614
rect 217222 660378 217306 660614
rect 217542 660378 250986 660614
rect 251222 660378 251306 660614
rect 251542 660378 284986 660614
rect 285222 660378 285306 660614
rect 285542 660378 318986 660614
rect 319222 660378 319306 660614
rect 319542 660378 352986 660614
rect 353222 660378 353306 660614
rect 353542 660378 386986 660614
rect 387222 660378 387306 660614
rect 387542 660378 420986 660614
rect 421222 660378 421306 660614
rect 421542 660378 454986 660614
rect 455222 660378 455306 660614
rect 455542 660378 488986 660614
rect 489222 660378 489306 660614
rect 489542 660378 522986 660614
rect 523222 660378 523306 660614
rect 523542 660378 556986 660614
rect 557222 660378 557306 660614
rect 557542 660378 588222 660614
rect 588458 660378 588542 660614
rect 588778 660378 592650 660614
rect -8726 660294 592650 660378
rect -8726 660058 -4854 660294
rect -4618 660058 -4534 660294
rect -4298 660058 12986 660294
rect 13222 660058 13306 660294
rect 13542 660058 46986 660294
rect 47222 660058 47306 660294
rect 47542 660058 80986 660294
rect 81222 660058 81306 660294
rect 81542 660058 114986 660294
rect 115222 660058 115306 660294
rect 115542 660058 148986 660294
rect 149222 660058 149306 660294
rect 149542 660058 182986 660294
rect 183222 660058 183306 660294
rect 183542 660058 216986 660294
rect 217222 660058 217306 660294
rect 217542 660058 250986 660294
rect 251222 660058 251306 660294
rect 251542 660058 284986 660294
rect 285222 660058 285306 660294
rect 285542 660058 318986 660294
rect 319222 660058 319306 660294
rect 319542 660058 352986 660294
rect 353222 660058 353306 660294
rect 353542 660058 386986 660294
rect 387222 660058 387306 660294
rect 387542 660058 420986 660294
rect 421222 660058 421306 660294
rect 421542 660058 454986 660294
rect 455222 660058 455306 660294
rect 455542 660058 488986 660294
rect 489222 660058 489306 660294
rect 489542 660058 522986 660294
rect 523222 660058 523306 660294
rect 523542 660058 556986 660294
rect 557222 660058 557306 660294
rect 557542 660058 588222 660294
rect 588458 660058 588542 660294
rect 588778 660058 592650 660294
rect -8726 660026 592650 660058
rect -8726 656894 592650 656926
rect -8726 656658 -3894 656894
rect -3658 656658 -3574 656894
rect -3338 656658 9266 656894
rect 9502 656658 9586 656894
rect 9822 656658 43266 656894
rect 43502 656658 43586 656894
rect 43822 656658 77266 656894
rect 77502 656658 77586 656894
rect 77822 656658 111266 656894
rect 111502 656658 111586 656894
rect 111822 656658 145266 656894
rect 145502 656658 145586 656894
rect 145822 656658 179266 656894
rect 179502 656658 179586 656894
rect 179822 656658 213266 656894
rect 213502 656658 213586 656894
rect 213822 656658 247266 656894
rect 247502 656658 247586 656894
rect 247822 656658 281266 656894
rect 281502 656658 281586 656894
rect 281822 656658 315266 656894
rect 315502 656658 315586 656894
rect 315822 656658 349266 656894
rect 349502 656658 349586 656894
rect 349822 656658 383266 656894
rect 383502 656658 383586 656894
rect 383822 656658 417266 656894
rect 417502 656658 417586 656894
rect 417822 656658 451266 656894
rect 451502 656658 451586 656894
rect 451822 656658 485266 656894
rect 485502 656658 485586 656894
rect 485822 656658 519266 656894
rect 519502 656658 519586 656894
rect 519822 656658 553266 656894
rect 553502 656658 553586 656894
rect 553822 656658 587262 656894
rect 587498 656658 587582 656894
rect 587818 656658 592650 656894
rect -8726 656574 592650 656658
rect -8726 656338 -3894 656574
rect -3658 656338 -3574 656574
rect -3338 656338 9266 656574
rect 9502 656338 9586 656574
rect 9822 656338 43266 656574
rect 43502 656338 43586 656574
rect 43822 656338 77266 656574
rect 77502 656338 77586 656574
rect 77822 656338 111266 656574
rect 111502 656338 111586 656574
rect 111822 656338 145266 656574
rect 145502 656338 145586 656574
rect 145822 656338 179266 656574
rect 179502 656338 179586 656574
rect 179822 656338 213266 656574
rect 213502 656338 213586 656574
rect 213822 656338 247266 656574
rect 247502 656338 247586 656574
rect 247822 656338 281266 656574
rect 281502 656338 281586 656574
rect 281822 656338 315266 656574
rect 315502 656338 315586 656574
rect 315822 656338 349266 656574
rect 349502 656338 349586 656574
rect 349822 656338 383266 656574
rect 383502 656338 383586 656574
rect 383822 656338 417266 656574
rect 417502 656338 417586 656574
rect 417822 656338 451266 656574
rect 451502 656338 451586 656574
rect 451822 656338 485266 656574
rect 485502 656338 485586 656574
rect 485822 656338 519266 656574
rect 519502 656338 519586 656574
rect 519822 656338 553266 656574
rect 553502 656338 553586 656574
rect 553822 656338 587262 656574
rect 587498 656338 587582 656574
rect 587818 656338 592650 656574
rect -8726 656306 592650 656338
rect -8726 653174 592650 653206
rect -8726 652938 -2934 653174
rect -2698 652938 -2614 653174
rect -2378 652938 5546 653174
rect 5782 652938 5866 653174
rect 6102 652938 39546 653174
rect 39782 652938 39866 653174
rect 40102 652938 73546 653174
rect 73782 652938 73866 653174
rect 74102 652938 107546 653174
rect 107782 652938 107866 653174
rect 108102 652938 141546 653174
rect 141782 652938 141866 653174
rect 142102 652938 175546 653174
rect 175782 652938 175866 653174
rect 176102 652938 209546 653174
rect 209782 652938 209866 653174
rect 210102 652938 243546 653174
rect 243782 652938 243866 653174
rect 244102 652938 277546 653174
rect 277782 652938 277866 653174
rect 278102 652938 311546 653174
rect 311782 652938 311866 653174
rect 312102 652938 345546 653174
rect 345782 652938 345866 653174
rect 346102 652938 379546 653174
rect 379782 652938 379866 653174
rect 380102 652938 413546 653174
rect 413782 652938 413866 653174
rect 414102 652938 447546 653174
rect 447782 652938 447866 653174
rect 448102 652938 481546 653174
rect 481782 652938 481866 653174
rect 482102 652938 515546 653174
rect 515782 652938 515866 653174
rect 516102 652938 549546 653174
rect 549782 652938 549866 653174
rect 550102 652938 586302 653174
rect 586538 652938 586622 653174
rect 586858 652938 592650 653174
rect -8726 652854 592650 652938
rect -8726 652618 -2934 652854
rect -2698 652618 -2614 652854
rect -2378 652618 5546 652854
rect 5782 652618 5866 652854
rect 6102 652618 39546 652854
rect 39782 652618 39866 652854
rect 40102 652618 73546 652854
rect 73782 652618 73866 652854
rect 74102 652618 107546 652854
rect 107782 652618 107866 652854
rect 108102 652618 141546 652854
rect 141782 652618 141866 652854
rect 142102 652618 175546 652854
rect 175782 652618 175866 652854
rect 176102 652618 209546 652854
rect 209782 652618 209866 652854
rect 210102 652618 243546 652854
rect 243782 652618 243866 652854
rect 244102 652618 277546 652854
rect 277782 652618 277866 652854
rect 278102 652618 311546 652854
rect 311782 652618 311866 652854
rect 312102 652618 345546 652854
rect 345782 652618 345866 652854
rect 346102 652618 379546 652854
rect 379782 652618 379866 652854
rect 380102 652618 413546 652854
rect 413782 652618 413866 652854
rect 414102 652618 447546 652854
rect 447782 652618 447866 652854
rect 448102 652618 481546 652854
rect 481782 652618 481866 652854
rect 482102 652618 515546 652854
rect 515782 652618 515866 652854
rect 516102 652618 549546 652854
rect 549782 652618 549866 652854
rect 550102 652618 586302 652854
rect 586538 652618 586622 652854
rect 586858 652618 592650 652854
rect -8726 652586 592650 652618
rect -8726 649454 592650 649486
rect -8726 649218 -1974 649454
rect -1738 649218 -1654 649454
rect -1418 649218 1826 649454
rect 2062 649218 2146 649454
rect 2382 649218 35826 649454
rect 36062 649218 36146 649454
rect 36382 649218 69826 649454
rect 70062 649218 70146 649454
rect 70382 649218 103826 649454
rect 104062 649218 104146 649454
rect 104382 649218 137826 649454
rect 138062 649218 138146 649454
rect 138382 649218 171826 649454
rect 172062 649218 172146 649454
rect 172382 649218 205826 649454
rect 206062 649218 206146 649454
rect 206382 649218 239826 649454
rect 240062 649218 240146 649454
rect 240382 649218 273826 649454
rect 274062 649218 274146 649454
rect 274382 649218 307826 649454
rect 308062 649218 308146 649454
rect 308382 649218 341826 649454
rect 342062 649218 342146 649454
rect 342382 649218 375826 649454
rect 376062 649218 376146 649454
rect 376382 649218 409826 649454
rect 410062 649218 410146 649454
rect 410382 649218 443826 649454
rect 444062 649218 444146 649454
rect 444382 649218 477826 649454
rect 478062 649218 478146 649454
rect 478382 649218 511826 649454
rect 512062 649218 512146 649454
rect 512382 649218 545826 649454
rect 546062 649218 546146 649454
rect 546382 649218 579826 649454
rect 580062 649218 580146 649454
rect 580382 649218 585342 649454
rect 585578 649218 585662 649454
rect 585898 649218 592650 649454
rect -8726 649134 592650 649218
rect -8726 648898 -1974 649134
rect -1738 648898 -1654 649134
rect -1418 648898 1826 649134
rect 2062 648898 2146 649134
rect 2382 648898 35826 649134
rect 36062 648898 36146 649134
rect 36382 648898 69826 649134
rect 70062 648898 70146 649134
rect 70382 648898 103826 649134
rect 104062 648898 104146 649134
rect 104382 648898 137826 649134
rect 138062 648898 138146 649134
rect 138382 648898 171826 649134
rect 172062 648898 172146 649134
rect 172382 648898 205826 649134
rect 206062 648898 206146 649134
rect 206382 648898 239826 649134
rect 240062 648898 240146 649134
rect 240382 648898 273826 649134
rect 274062 648898 274146 649134
rect 274382 648898 307826 649134
rect 308062 648898 308146 649134
rect 308382 648898 341826 649134
rect 342062 648898 342146 649134
rect 342382 648898 375826 649134
rect 376062 648898 376146 649134
rect 376382 648898 409826 649134
rect 410062 648898 410146 649134
rect 410382 648898 443826 649134
rect 444062 648898 444146 649134
rect 444382 648898 477826 649134
rect 478062 648898 478146 649134
rect 478382 648898 511826 649134
rect 512062 648898 512146 649134
rect 512382 648898 545826 649134
rect 546062 648898 546146 649134
rect 546382 648898 579826 649134
rect 580062 648898 580146 649134
rect 580382 648898 585342 649134
rect 585578 648898 585662 649134
rect 585898 648898 592650 649134
rect -8726 648866 592650 648898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 61866 641494
rect 62102 641258 62186 641494
rect 62422 641258 95866 641494
rect 96102 641258 96186 641494
rect 96422 641258 129866 641494
rect 130102 641258 130186 641494
rect 130422 641258 163866 641494
rect 164102 641258 164186 641494
rect 164422 641258 197866 641494
rect 198102 641258 198186 641494
rect 198422 641258 231866 641494
rect 232102 641258 232186 641494
rect 232422 641258 265866 641494
rect 266102 641258 266186 641494
rect 266422 641258 299866 641494
rect 300102 641258 300186 641494
rect 300422 641258 333866 641494
rect 334102 641258 334186 641494
rect 334422 641258 367866 641494
rect 368102 641258 368186 641494
rect 368422 641258 401866 641494
rect 402102 641258 402186 641494
rect 402422 641258 435866 641494
rect 436102 641258 436186 641494
rect 436422 641258 469866 641494
rect 470102 641258 470186 641494
rect 470422 641258 503866 641494
rect 504102 641258 504186 641494
rect 504422 641258 537866 641494
rect 538102 641258 538186 641494
rect 538422 641258 571866 641494
rect 572102 641258 572186 641494
rect 572422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 61866 641174
rect 62102 640938 62186 641174
rect 62422 640938 95866 641174
rect 96102 640938 96186 641174
rect 96422 640938 129866 641174
rect 130102 640938 130186 641174
rect 130422 640938 163866 641174
rect 164102 640938 164186 641174
rect 164422 640938 197866 641174
rect 198102 640938 198186 641174
rect 198422 640938 231866 641174
rect 232102 640938 232186 641174
rect 232422 640938 265866 641174
rect 266102 640938 266186 641174
rect 266422 640938 299866 641174
rect 300102 640938 300186 641174
rect 300422 640938 333866 641174
rect 334102 640938 334186 641174
rect 334422 640938 367866 641174
rect 368102 640938 368186 641174
rect 368422 640938 401866 641174
rect 402102 640938 402186 641174
rect 402422 640938 435866 641174
rect 436102 640938 436186 641174
rect 436422 640938 469866 641174
rect 470102 640938 470186 641174
rect 470422 640938 503866 641174
rect 504102 640938 504186 641174
rect 504422 640938 537866 641174
rect 538102 640938 538186 641174
rect 538422 640938 571866 641174
rect 572102 640938 572186 641174
rect 572422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 58146 637774
rect 58382 637538 58466 637774
rect 58702 637538 92146 637774
rect 92382 637538 92466 637774
rect 92702 637538 126146 637774
rect 126382 637538 126466 637774
rect 126702 637538 160146 637774
rect 160382 637538 160466 637774
rect 160702 637538 194146 637774
rect 194382 637538 194466 637774
rect 194702 637538 228146 637774
rect 228382 637538 228466 637774
rect 228702 637538 262146 637774
rect 262382 637538 262466 637774
rect 262702 637538 296146 637774
rect 296382 637538 296466 637774
rect 296702 637538 330146 637774
rect 330382 637538 330466 637774
rect 330702 637538 364146 637774
rect 364382 637538 364466 637774
rect 364702 637538 398146 637774
rect 398382 637538 398466 637774
rect 398702 637538 432146 637774
rect 432382 637538 432466 637774
rect 432702 637538 466146 637774
rect 466382 637538 466466 637774
rect 466702 637538 500146 637774
rect 500382 637538 500466 637774
rect 500702 637538 534146 637774
rect 534382 637538 534466 637774
rect 534702 637538 568146 637774
rect 568382 637538 568466 637774
rect 568702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 58146 637454
rect 58382 637218 58466 637454
rect 58702 637218 92146 637454
rect 92382 637218 92466 637454
rect 92702 637218 126146 637454
rect 126382 637218 126466 637454
rect 126702 637218 160146 637454
rect 160382 637218 160466 637454
rect 160702 637218 194146 637454
rect 194382 637218 194466 637454
rect 194702 637218 228146 637454
rect 228382 637218 228466 637454
rect 228702 637218 262146 637454
rect 262382 637218 262466 637454
rect 262702 637218 296146 637454
rect 296382 637218 296466 637454
rect 296702 637218 330146 637454
rect 330382 637218 330466 637454
rect 330702 637218 364146 637454
rect 364382 637218 364466 637454
rect 364702 637218 398146 637454
rect 398382 637218 398466 637454
rect 398702 637218 432146 637454
rect 432382 637218 432466 637454
rect 432702 637218 466146 637454
rect 466382 637218 466466 637454
rect 466702 637218 500146 637454
rect 500382 637218 500466 637454
rect 500702 637218 534146 637454
rect 534382 637218 534466 637454
rect 534702 637218 568146 637454
rect 568382 637218 568466 637454
rect 568702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 54426 634054
rect 54662 633818 54746 634054
rect 54982 633818 88426 634054
rect 88662 633818 88746 634054
rect 88982 633818 122426 634054
rect 122662 633818 122746 634054
rect 122982 633818 156426 634054
rect 156662 633818 156746 634054
rect 156982 633818 190426 634054
rect 190662 633818 190746 634054
rect 190982 633818 224426 634054
rect 224662 633818 224746 634054
rect 224982 633818 258426 634054
rect 258662 633818 258746 634054
rect 258982 633818 292426 634054
rect 292662 633818 292746 634054
rect 292982 633818 326426 634054
rect 326662 633818 326746 634054
rect 326982 633818 360426 634054
rect 360662 633818 360746 634054
rect 360982 633818 394426 634054
rect 394662 633818 394746 634054
rect 394982 633818 428426 634054
rect 428662 633818 428746 634054
rect 428982 633818 462426 634054
rect 462662 633818 462746 634054
rect 462982 633818 496426 634054
rect 496662 633818 496746 634054
rect 496982 633818 530426 634054
rect 530662 633818 530746 634054
rect 530982 633818 564426 634054
rect 564662 633818 564746 634054
rect 564982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 54426 633734
rect 54662 633498 54746 633734
rect 54982 633498 88426 633734
rect 88662 633498 88746 633734
rect 88982 633498 122426 633734
rect 122662 633498 122746 633734
rect 122982 633498 156426 633734
rect 156662 633498 156746 633734
rect 156982 633498 190426 633734
rect 190662 633498 190746 633734
rect 190982 633498 224426 633734
rect 224662 633498 224746 633734
rect 224982 633498 258426 633734
rect 258662 633498 258746 633734
rect 258982 633498 292426 633734
rect 292662 633498 292746 633734
rect 292982 633498 326426 633734
rect 326662 633498 326746 633734
rect 326982 633498 360426 633734
rect 360662 633498 360746 633734
rect 360982 633498 394426 633734
rect 394662 633498 394746 633734
rect 394982 633498 428426 633734
rect 428662 633498 428746 633734
rect 428982 633498 462426 633734
rect 462662 633498 462746 633734
rect 462982 633498 496426 633734
rect 496662 633498 496746 633734
rect 496982 633498 530426 633734
rect 530662 633498 530746 633734
rect 530982 633498 564426 633734
rect 564662 633498 564746 633734
rect 564982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 50706 630334
rect 50942 630098 51026 630334
rect 51262 630098 84706 630334
rect 84942 630098 85026 630334
rect 85262 630098 118706 630334
rect 118942 630098 119026 630334
rect 119262 630098 152706 630334
rect 152942 630098 153026 630334
rect 153262 630098 186706 630334
rect 186942 630098 187026 630334
rect 187262 630098 220706 630334
rect 220942 630098 221026 630334
rect 221262 630098 254706 630334
rect 254942 630098 255026 630334
rect 255262 630098 288706 630334
rect 288942 630098 289026 630334
rect 289262 630098 322706 630334
rect 322942 630098 323026 630334
rect 323262 630098 356706 630334
rect 356942 630098 357026 630334
rect 357262 630098 390706 630334
rect 390942 630098 391026 630334
rect 391262 630098 424706 630334
rect 424942 630098 425026 630334
rect 425262 630098 458706 630334
rect 458942 630098 459026 630334
rect 459262 630098 492706 630334
rect 492942 630098 493026 630334
rect 493262 630098 526706 630334
rect 526942 630098 527026 630334
rect 527262 630098 560706 630334
rect 560942 630098 561026 630334
rect 561262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 50706 630014
rect 50942 629778 51026 630014
rect 51262 629778 84706 630014
rect 84942 629778 85026 630014
rect 85262 629778 118706 630014
rect 118942 629778 119026 630014
rect 119262 629778 152706 630014
rect 152942 629778 153026 630014
rect 153262 629778 186706 630014
rect 186942 629778 187026 630014
rect 187262 629778 220706 630014
rect 220942 629778 221026 630014
rect 221262 629778 254706 630014
rect 254942 629778 255026 630014
rect 255262 629778 288706 630014
rect 288942 629778 289026 630014
rect 289262 629778 322706 630014
rect 322942 629778 323026 630014
rect 323262 629778 356706 630014
rect 356942 629778 357026 630014
rect 357262 629778 390706 630014
rect 390942 629778 391026 630014
rect 391262 629778 424706 630014
rect 424942 629778 425026 630014
rect 425262 629778 458706 630014
rect 458942 629778 459026 630014
rect 459262 629778 492706 630014
rect 492942 629778 493026 630014
rect 493262 629778 526706 630014
rect 526942 629778 527026 630014
rect 527262 629778 560706 630014
rect 560942 629778 561026 630014
rect 561262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 46986 626614
rect 47222 626378 47306 626614
rect 47542 626378 80986 626614
rect 81222 626378 81306 626614
rect 81542 626378 114986 626614
rect 115222 626378 115306 626614
rect 115542 626378 148986 626614
rect 149222 626378 149306 626614
rect 149542 626378 182986 626614
rect 183222 626378 183306 626614
rect 183542 626378 216986 626614
rect 217222 626378 217306 626614
rect 217542 626378 250986 626614
rect 251222 626378 251306 626614
rect 251542 626378 284986 626614
rect 285222 626378 285306 626614
rect 285542 626378 318986 626614
rect 319222 626378 319306 626614
rect 319542 626378 352986 626614
rect 353222 626378 353306 626614
rect 353542 626378 386986 626614
rect 387222 626378 387306 626614
rect 387542 626378 420986 626614
rect 421222 626378 421306 626614
rect 421542 626378 454986 626614
rect 455222 626378 455306 626614
rect 455542 626378 488986 626614
rect 489222 626378 489306 626614
rect 489542 626378 522986 626614
rect 523222 626378 523306 626614
rect 523542 626378 556986 626614
rect 557222 626378 557306 626614
rect 557542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 46986 626294
rect 47222 626058 47306 626294
rect 47542 626058 80986 626294
rect 81222 626058 81306 626294
rect 81542 626058 114986 626294
rect 115222 626058 115306 626294
rect 115542 626058 148986 626294
rect 149222 626058 149306 626294
rect 149542 626058 182986 626294
rect 183222 626058 183306 626294
rect 183542 626058 216986 626294
rect 217222 626058 217306 626294
rect 217542 626058 250986 626294
rect 251222 626058 251306 626294
rect 251542 626058 284986 626294
rect 285222 626058 285306 626294
rect 285542 626058 318986 626294
rect 319222 626058 319306 626294
rect 319542 626058 352986 626294
rect 353222 626058 353306 626294
rect 353542 626058 386986 626294
rect 387222 626058 387306 626294
rect 387542 626058 420986 626294
rect 421222 626058 421306 626294
rect 421542 626058 454986 626294
rect 455222 626058 455306 626294
rect 455542 626058 488986 626294
rect 489222 626058 489306 626294
rect 489542 626058 522986 626294
rect 523222 626058 523306 626294
rect 523542 626058 556986 626294
rect 557222 626058 557306 626294
rect 557542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 43266 622894
rect 43502 622658 43586 622894
rect 43822 622658 77266 622894
rect 77502 622658 77586 622894
rect 77822 622658 111266 622894
rect 111502 622658 111586 622894
rect 111822 622658 145266 622894
rect 145502 622658 145586 622894
rect 145822 622658 179266 622894
rect 179502 622658 179586 622894
rect 179822 622658 213266 622894
rect 213502 622658 213586 622894
rect 213822 622658 247266 622894
rect 247502 622658 247586 622894
rect 247822 622658 281266 622894
rect 281502 622658 281586 622894
rect 281822 622658 315266 622894
rect 315502 622658 315586 622894
rect 315822 622658 349266 622894
rect 349502 622658 349586 622894
rect 349822 622658 383266 622894
rect 383502 622658 383586 622894
rect 383822 622658 417266 622894
rect 417502 622658 417586 622894
rect 417822 622658 451266 622894
rect 451502 622658 451586 622894
rect 451822 622658 485266 622894
rect 485502 622658 485586 622894
rect 485822 622658 519266 622894
rect 519502 622658 519586 622894
rect 519822 622658 553266 622894
rect 553502 622658 553586 622894
rect 553822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 43266 622574
rect 43502 622338 43586 622574
rect 43822 622338 77266 622574
rect 77502 622338 77586 622574
rect 77822 622338 111266 622574
rect 111502 622338 111586 622574
rect 111822 622338 145266 622574
rect 145502 622338 145586 622574
rect 145822 622338 179266 622574
rect 179502 622338 179586 622574
rect 179822 622338 213266 622574
rect 213502 622338 213586 622574
rect 213822 622338 247266 622574
rect 247502 622338 247586 622574
rect 247822 622338 281266 622574
rect 281502 622338 281586 622574
rect 281822 622338 315266 622574
rect 315502 622338 315586 622574
rect 315822 622338 349266 622574
rect 349502 622338 349586 622574
rect 349822 622338 383266 622574
rect 383502 622338 383586 622574
rect 383822 622338 417266 622574
rect 417502 622338 417586 622574
rect 417822 622338 451266 622574
rect 451502 622338 451586 622574
rect 451822 622338 485266 622574
rect 485502 622338 485586 622574
rect 485822 622338 519266 622574
rect 519502 622338 519586 622574
rect 519822 622338 553266 622574
rect 553502 622338 553586 622574
rect 553822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39546 619174
rect 39782 618938 39866 619174
rect 40102 618938 73546 619174
rect 73782 618938 73866 619174
rect 74102 618938 107546 619174
rect 107782 618938 107866 619174
rect 108102 618938 141546 619174
rect 141782 618938 141866 619174
rect 142102 618938 175546 619174
rect 175782 618938 175866 619174
rect 176102 618938 209546 619174
rect 209782 618938 209866 619174
rect 210102 618938 243546 619174
rect 243782 618938 243866 619174
rect 244102 618938 277546 619174
rect 277782 618938 277866 619174
rect 278102 618938 311546 619174
rect 311782 618938 311866 619174
rect 312102 618938 345546 619174
rect 345782 618938 345866 619174
rect 346102 618938 379546 619174
rect 379782 618938 379866 619174
rect 380102 618938 413546 619174
rect 413782 618938 413866 619174
rect 414102 618938 447546 619174
rect 447782 618938 447866 619174
rect 448102 618938 481546 619174
rect 481782 618938 481866 619174
rect 482102 618938 515546 619174
rect 515782 618938 515866 619174
rect 516102 618938 549546 619174
rect 549782 618938 549866 619174
rect 550102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39546 618854
rect 39782 618618 39866 618854
rect 40102 618618 73546 618854
rect 73782 618618 73866 618854
rect 74102 618618 107546 618854
rect 107782 618618 107866 618854
rect 108102 618618 141546 618854
rect 141782 618618 141866 618854
rect 142102 618618 175546 618854
rect 175782 618618 175866 618854
rect 176102 618618 209546 618854
rect 209782 618618 209866 618854
rect 210102 618618 243546 618854
rect 243782 618618 243866 618854
rect 244102 618618 277546 618854
rect 277782 618618 277866 618854
rect 278102 618618 311546 618854
rect 311782 618618 311866 618854
rect 312102 618618 345546 618854
rect 345782 618618 345866 618854
rect 346102 618618 379546 618854
rect 379782 618618 379866 618854
rect 380102 618618 413546 618854
rect 413782 618618 413866 618854
rect 414102 618618 447546 618854
rect 447782 618618 447866 618854
rect 448102 618618 481546 618854
rect 481782 618618 481866 618854
rect 482102 618618 515546 618854
rect 515782 618618 515866 618854
rect 516102 618618 549546 618854
rect 549782 618618 549866 618854
rect 550102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 35826 615454
rect 36062 615218 36146 615454
rect 36382 615218 69826 615454
rect 70062 615218 70146 615454
rect 70382 615218 103826 615454
rect 104062 615218 104146 615454
rect 104382 615218 137826 615454
rect 138062 615218 138146 615454
rect 138382 615218 171826 615454
rect 172062 615218 172146 615454
rect 172382 615218 205826 615454
rect 206062 615218 206146 615454
rect 206382 615218 239826 615454
rect 240062 615218 240146 615454
rect 240382 615218 273826 615454
rect 274062 615218 274146 615454
rect 274382 615218 307826 615454
rect 308062 615218 308146 615454
rect 308382 615218 341826 615454
rect 342062 615218 342146 615454
rect 342382 615218 375826 615454
rect 376062 615218 376146 615454
rect 376382 615218 409826 615454
rect 410062 615218 410146 615454
rect 410382 615218 443826 615454
rect 444062 615218 444146 615454
rect 444382 615218 477826 615454
rect 478062 615218 478146 615454
rect 478382 615218 511826 615454
rect 512062 615218 512146 615454
rect 512382 615218 545826 615454
rect 546062 615218 546146 615454
rect 546382 615218 579826 615454
rect 580062 615218 580146 615454
rect 580382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 35826 615134
rect 36062 614898 36146 615134
rect 36382 614898 69826 615134
rect 70062 614898 70146 615134
rect 70382 614898 103826 615134
rect 104062 614898 104146 615134
rect 104382 614898 137826 615134
rect 138062 614898 138146 615134
rect 138382 614898 171826 615134
rect 172062 614898 172146 615134
rect 172382 614898 205826 615134
rect 206062 614898 206146 615134
rect 206382 614898 239826 615134
rect 240062 614898 240146 615134
rect 240382 614898 273826 615134
rect 274062 614898 274146 615134
rect 274382 614898 307826 615134
rect 308062 614898 308146 615134
rect 308382 614898 341826 615134
rect 342062 614898 342146 615134
rect 342382 614898 375826 615134
rect 376062 614898 376146 615134
rect 376382 614898 409826 615134
rect 410062 614898 410146 615134
rect 410382 614898 443826 615134
rect 444062 614898 444146 615134
rect 444382 614898 477826 615134
rect 478062 614898 478146 615134
rect 478382 614898 511826 615134
rect 512062 614898 512146 615134
rect 512382 614898 545826 615134
rect 546062 614898 546146 615134
rect 546382 614898 579826 615134
rect 580062 614898 580146 615134
rect 580382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 607494 592650 607526
rect -8726 607258 -8694 607494
rect -8458 607258 -8374 607494
rect -8138 607258 27866 607494
rect 28102 607258 28186 607494
rect 28422 607258 61866 607494
rect 62102 607258 62186 607494
rect 62422 607258 95866 607494
rect 96102 607258 96186 607494
rect 96422 607258 129866 607494
rect 130102 607258 130186 607494
rect 130422 607258 163866 607494
rect 164102 607258 164186 607494
rect 164422 607258 197866 607494
rect 198102 607258 198186 607494
rect 198422 607258 231866 607494
rect 232102 607258 232186 607494
rect 232422 607258 265866 607494
rect 266102 607258 266186 607494
rect 266422 607258 299866 607494
rect 300102 607258 300186 607494
rect 300422 607258 333866 607494
rect 334102 607258 334186 607494
rect 334422 607258 367866 607494
rect 368102 607258 368186 607494
rect 368422 607258 401866 607494
rect 402102 607258 402186 607494
rect 402422 607258 435866 607494
rect 436102 607258 436186 607494
rect 436422 607258 469866 607494
rect 470102 607258 470186 607494
rect 470422 607258 503866 607494
rect 504102 607258 504186 607494
rect 504422 607258 537866 607494
rect 538102 607258 538186 607494
rect 538422 607258 571866 607494
rect 572102 607258 572186 607494
rect 572422 607258 592062 607494
rect 592298 607258 592382 607494
rect 592618 607258 592650 607494
rect -8726 607174 592650 607258
rect -8726 606938 -8694 607174
rect -8458 606938 -8374 607174
rect -8138 606938 27866 607174
rect 28102 606938 28186 607174
rect 28422 606938 61866 607174
rect 62102 606938 62186 607174
rect 62422 606938 95866 607174
rect 96102 606938 96186 607174
rect 96422 606938 129866 607174
rect 130102 606938 130186 607174
rect 130422 606938 163866 607174
rect 164102 606938 164186 607174
rect 164422 606938 197866 607174
rect 198102 606938 198186 607174
rect 198422 606938 231866 607174
rect 232102 606938 232186 607174
rect 232422 606938 265866 607174
rect 266102 606938 266186 607174
rect 266422 606938 299866 607174
rect 300102 606938 300186 607174
rect 300422 606938 333866 607174
rect 334102 606938 334186 607174
rect 334422 606938 367866 607174
rect 368102 606938 368186 607174
rect 368422 606938 401866 607174
rect 402102 606938 402186 607174
rect 402422 606938 435866 607174
rect 436102 606938 436186 607174
rect 436422 606938 469866 607174
rect 470102 606938 470186 607174
rect 470422 606938 503866 607174
rect 504102 606938 504186 607174
rect 504422 606938 537866 607174
rect 538102 606938 538186 607174
rect 538422 606938 571866 607174
rect 572102 606938 572186 607174
rect 572422 606938 592062 607174
rect 592298 606938 592382 607174
rect 592618 606938 592650 607174
rect -8726 606906 592650 606938
rect -8726 603774 592650 603806
rect -8726 603538 -7734 603774
rect -7498 603538 -7414 603774
rect -7178 603538 24146 603774
rect 24382 603538 24466 603774
rect 24702 603538 58146 603774
rect 58382 603538 58466 603774
rect 58702 603538 92146 603774
rect 92382 603538 92466 603774
rect 92702 603538 126146 603774
rect 126382 603538 126466 603774
rect 126702 603538 160146 603774
rect 160382 603538 160466 603774
rect 160702 603538 194146 603774
rect 194382 603538 194466 603774
rect 194702 603538 228146 603774
rect 228382 603538 228466 603774
rect 228702 603538 262146 603774
rect 262382 603538 262466 603774
rect 262702 603538 296146 603774
rect 296382 603538 296466 603774
rect 296702 603538 330146 603774
rect 330382 603538 330466 603774
rect 330702 603538 364146 603774
rect 364382 603538 364466 603774
rect 364702 603538 398146 603774
rect 398382 603538 398466 603774
rect 398702 603538 432146 603774
rect 432382 603538 432466 603774
rect 432702 603538 466146 603774
rect 466382 603538 466466 603774
rect 466702 603538 500146 603774
rect 500382 603538 500466 603774
rect 500702 603538 534146 603774
rect 534382 603538 534466 603774
rect 534702 603538 568146 603774
rect 568382 603538 568466 603774
rect 568702 603538 591102 603774
rect 591338 603538 591422 603774
rect 591658 603538 592650 603774
rect -8726 603454 592650 603538
rect -8726 603218 -7734 603454
rect -7498 603218 -7414 603454
rect -7178 603218 24146 603454
rect 24382 603218 24466 603454
rect 24702 603218 58146 603454
rect 58382 603218 58466 603454
rect 58702 603218 92146 603454
rect 92382 603218 92466 603454
rect 92702 603218 126146 603454
rect 126382 603218 126466 603454
rect 126702 603218 160146 603454
rect 160382 603218 160466 603454
rect 160702 603218 194146 603454
rect 194382 603218 194466 603454
rect 194702 603218 228146 603454
rect 228382 603218 228466 603454
rect 228702 603218 262146 603454
rect 262382 603218 262466 603454
rect 262702 603218 296146 603454
rect 296382 603218 296466 603454
rect 296702 603218 330146 603454
rect 330382 603218 330466 603454
rect 330702 603218 364146 603454
rect 364382 603218 364466 603454
rect 364702 603218 398146 603454
rect 398382 603218 398466 603454
rect 398702 603218 432146 603454
rect 432382 603218 432466 603454
rect 432702 603218 466146 603454
rect 466382 603218 466466 603454
rect 466702 603218 500146 603454
rect 500382 603218 500466 603454
rect 500702 603218 534146 603454
rect 534382 603218 534466 603454
rect 534702 603218 568146 603454
rect 568382 603218 568466 603454
rect 568702 603218 591102 603454
rect 591338 603218 591422 603454
rect 591658 603218 592650 603454
rect -8726 603186 592650 603218
rect -8726 600054 592650 600086
rect -8726 599818 -6774 600054
rect -6538 599818 -6454 600054
rect -6218 599818 20426 600054
rect 20662 599818 20746 600054
rect 20982 599818 54426 600054
rect 54662 599818 54746 600054
rect 54982 599818 88426 600054
rect 88662 599818 88746 600054
rect 88982 599818 122426 600054
rect 122662 599818 122746 600054
rect 122982 599818 156426 600054
rect 156662 599818 156746 600054
rect 156982 599818 190426 600054
rect 190662 599818 190746 600054
rect 190982 599818 224426 600054
rect 224662 599818 224746 600054
rect 224982 599818 258426 600054
rect 258662 599818 258746 600054
rect 258982 599818 292426 600054
rect 292662 599818 292746 600054
rect 292982 599818 326426 600054
rect 326662 599818 326746 600054
rect 326982 599818 360426 600054
rect 360662 599818 360746 600054
rect 360982 599818 394426 600054
rect 394662 599818 394746 600054
rect 394982 599818 428426 600054
rect 428662 599818 428746 600054
rect 428982 599818 462426 600054
rect 462662 599818 462746 600054
rect 462982 599818 496426 600054
rect 496662 599818 496746 600054
rect 496982 599818 530426 600054
rect 530662 599818 530746 600054
rect 530982 599818 564426 600054
rect 564662 599818 564746 600054
rect 564982 599818 590142 600054
rect 590378 599818 590462 600054
rect 590698 599818 592650 600054
rect -8726 599734 592650 599818
rect -8726 599498 -6774 599734
rect -6538 599498 -6454 599734
rect -6218 599498 20426 599734
rect 20662 599498 20746 599734
rect 20982 599498 54426 599734
rect 54662 599498 54746 599734
rect 54982 599498 88426 599734
rect 88662 599498 88746 599734
rect 88982 599498 122426 599734
rect 122662 599498 122746 599734
rect 122982 599498 156426 599734
rect 156662 599498 156746 599734
rect 156982 599498 190426 599734
rect 190662 599498 190746 599734
rect 190982 599498 224426 599734
rect 224662 599498 224746 599734
rect 224982 599498 258426 599734
rect 258662 599498 258746 599734
rect 258982 599498 292426 599734
rect 292662 599498 292746 599734
rect 292982 599498 326426 599734
rect 326662 599498 326746 599734
rect 326982 599498 360426 599734
rect 360662 599498 360746 599734
rect 360982 599498 394426 599734
rect 394662 599498 394746 599734
rect 394982 599498 428426 599734
rect 428662 599498 428746 599734
rect 428982 599498 462426 599734
rect 462662 599498 462746 599734
rect 462982 599498 496426 599734
rect 496662 599498 496746 599734
rect 496982 599498 530426 599734
rect 530662 599498 530746 599734
rect 530982 599498 564426 599734
rect 564662 599498 564746 599734
rect 564982 599498 590142 599734
rect 590378 599498 590462 599734
rect 590698 599498 592650 599734
rect -8726 599466 592650 599498
rect -8726 596334 592650 596366
rect -8726 596098 -5814 596334
rect -5578 596098 -5494 596334
rect -5258 596098 16706 596334
rect 16942 596098 17026 596334
rect 17262 596098 50706 596334
rect 50942 596098 51026 596334
rect 51262 596098 84706 596334
rect 84942 596098 85026 596334
rect 85262 596098 118706 596334
rect 118942 596098 119026 596334
rect 119262 596098 152706 596334
rect 152942 596098 153026 596334
rect 153262 596098 186706 596334
rect 186942 596098 187026 596334
rect 187262 596098 220706 596334
rect 220942 596098 221026 596334
rect 221262 596098 254706 596334
rect 254942 596098 255026 596334
rect 255262 596098 288706 596334
rect 288942 596098 289026 596334
rect 289262 596098 322706 596334
rect 322942 596098 323026 596334
rect 323262 596098 356706 596334
rect 356942 596098 357026 596334
rect 357262 596098 390706 596334
rect 390942 596098 391026 596334
rect 391262 596098 424706 596334
rect 424942 596098 425026 596334
rect 425262 596098 458706 596334
rect 458942 596098 459026 596334
rect 459262 596098 492706 596334
rect 492942 596098 493026 596334
rect 493262 596098 526706 596334
rect 526942 596098 527026 596334
rect 527262 596098 560706 596334
rect 560942 596098 561026 596334
rect 561262 596098 589182 596334
rect 589418 596098 589502 596334
rect 589738 596098 592650 596334
rect -8726 596014 592650 596098
rect -8726 595778 -5814 596014
rect -5578 595778 -5494 596014
rect -5258 595778 16706 596014
rect 16942 595778 17026 596014
rect 17262 595778 50706 596014
rect 50942 595778 51026 596014
rect 51262 595778 84706 596014
rect 84942 595778 85026 596014
rect 85262 595778 118706 596014
rect 118942 595778 119026 596014
rect 119262 595778 152706 596014
rect 152942 595778 153026 596014
rect 153262 595778 186706 596014
rect 186942 595778 187026 596014
rect 187262 595778 220706 596014
rect 220942 595778 221026 596014
rect 221262 595778 254706 596014
rect 254942 595778 255026 596014
rect 255262 595778 288706 596014
rect 288942 595778 289026 596014
rect 289262 595778 322706 596014
rect 322942 595778 323026 596014
rect 323262 595778 356706 596014
rect 356942 595778 357026 596014
rect 357262 595778 390706 596014
rect 390942 595778 391026 596014
rect 391262 595778 424706 596014
rect 424942 595778 425026 596014
rect 425262 595778 458706 596014
rect 458942 595778 459026 596014
rect 459262 595778 492706 596014
rect 492942 595778 493026 596014
rect 493262 595778 526706 596014
rect 526942 595778 527026 596014
rect 527262 595778 560706 596014
rect 560942 595778 561026 596014
rect 561262 595778 589182 596014
rect 589418 595778 589502 596014
rect 589738 595778 592650 596014
rect -8726 595746 592650 595778
rect -8726 592614 592650 592646
rect -8726 592378 -4854 592614
rect -4618 592378 -4534 592614
rect -4298 592378 12986 592614
rect 13222 592378 13306 592614
rect 13542 592378 46986 592614
rect 47222 592378 47306 592614
rect 47542 592378 80986 592614
rect 81222 592378 81306 592614
rect 81542 592378 114986 592614
rect 115222 592378 115306 592614
rect 115542 592378 148986 592614
rect 149222 592378 149306 592614
rect 149542 592378 182986 592614
rect 183222 592378 183306 592614
rect 183542 592378 216986 592614
rect 217222 592378 217306 592614
rect 217542 592378 250986 592614
rect 251222 592378 251306 592614
rect 251542 592378 284986 592614
rect 285222 592378 285306 592614
rect 285542 592378 318986 592614
rect 319222 592378 319306 592614
rect 319542 592378 352986 592614
rect 353222 592378 353306 592614
rect 353542 592378 386986 592614
rect 387222 592378 387306 592614
rect 387542 592378 420986 592614
rect 421222 592378 421306 592614
rect 421542 592378 454986 592614
rect 455222 592378 455306 592614
rect 455542 592378 488986 592614
rect 489222 592378 489306 592614
rect 489542 592378 522986 592614
rect 523222 592378 523306 592614
rect 523542 592378 556986 592614
rect 557222 592378 557306 592614
rect 557542 592378 588222 592614
rect 588458 592378 588542 592614
rect 588778 592378 592650 592614
rect -8726 592294 592650 592378
rect -8726 592058 -4854 592294
rect -4618 592058 -4534 592294
rect -4298 592058 12986 592294
rect 13222 592058 13306 592294
rect 13542 592058 46986 592294
rect 47222 592058 47306 592294
rect 47542 592058 80986 592294
rect 81222 592058 81306 592294
rect 81542 592058 114986 592294
rect 115222 592058 115306 592294
rect 115542 592058 148986 592294
rect 149222 592058 149306 592294
rect 149542 592058 182986 592294
rect 183222 592058 183306 592294
rect 183542 592058 216986 592294
rect 217222 592058 217306 592294
rect 217542 592058 250986 592294
rect 251222 592058 251306 592294
rect 251542 592058 284986 592294
rect 285222 592058 285306 592294
rect 285542 592058 318986 592294
rect 319222 592058 319306 592294
rect 319542 592058 352986 592294
rect 353222 592058 353306 592294
rect 353542 592058 386986 592294
rect 387222 592058 387306 592294
rect 387542 592058 420986 592294
rect 421222 592058 421306 592294
rect 421542 592058 454986 592294
rect 455222 592058 455306 592294
rect 455542 592058 488986 592294
rect 489222 592058 489306 592294
rect 489542 592058 522986 592294
rect 523222 592058 523306 592294
rect 523542 592058 556986 592294
rect 557222 592058 557306 592294
rect 557542 592058 588222 592294
rect 588458 592058 588542 592294
rect 588778 592058 592650 592294
rect -8726 592026 592650 592058
rect -8726 588894 592650 588926
rect -8726 588658 -3894 588894
rect -3658 588658 -3574 588894
rect -3338 588658 9266 588894
rect 9502 588658 9586 588894
rect 9822 588658 43266 588894
rect 43502 588658 43586 588894
rect 43822 588658 77266 588894
rect 77502 588658 77586 588894
rect 77822 588658 111266 588894
rect 111502 588658 111586 588894
rect 111822 588658 145266 588894
rect 145502 588658 145586 588894
rect 145822 588658 179266 588894
rect 179502 588658 179586 588894
rect 179822 588658 213266 588894
rect 213502 588658 213586 588894
rect 213822 588658 247266 588894
rect 247502 588658 247586 588894
rect 247822 588658 281266 588894
rect 281502 588658 281586 588894
rect 281822 588658 315266 588894
rect 315502 588658 315586 588894
rect 315822 588658 349266 588894
rect 349502 588658 349586 588894
rect 349822 588658 383266 588894
rect 383502 588658 383586 588894
rect 383822 588658 417266 588894
rect 417502 588658 417586 588894
rect 417822 588658 451266 588894
rect 451502 588658 451586 588894
rect 451822 588658 485266 588894
rect 485502 588658 485586 588894
rect 485822 588658 519266 588894
rect 519502 588658 519586 588894
rect 519822 588658 553266 588894
rect 553502 588658 553586 588894
rect 553822 588658 587262 588894
rect 587498 588658 587582 588894
rect 587818 588658 592650 588894
rect -8726 588574 592650 588658
rect -8726 588338 -3894 588574
rect -3658 588338 -3574 588574
rect -3338 588338 9266 588574
rect 9502 588338 9586 588574
rect 9822 588338 43266 588574
rect 43502 588338 43586 588574
rect 43822 588338 77266 588574
rect 77502 588338 77586 588574
rect 77822 588338 111266 588574
rect 111502 588338 111586 588574
rect 111822 588338 145266 588574
rect 145502 588338 145586 588574
rect 145822 588338 179266 588574
rect 179502 588338 179586 588574
rect 179822 588338 213266 588574
rect 213502 588338 213586 588574
rect 213822 588338 247266 588574
rect 247502 588338 247586 588574
rect 247822 588338 281266 588574
rect 281502 588338 281586 588574
rect 281822 588338 315266 588574
rect 315502 588338 315586 588574
rect 315822 588338 349266 588574
rect 349502 588338 349586 588574
rect 349822 588338 383266 588574
rect 383502 588338 383586 588574
rect 383822 588338 417266 588574
rect 417502 588338 417586 588574
rect 417822 588338 451266 588574
rect 451502 588338 451586 588574
rect 451822 588338 485266 588574
rect 485502 588338 485586 588574
rect 485822 588338 519266 588574
rect 519502 588338 519586 588574
rect 519822 588338 553266 588574
rect 553502 588338 553586 588574
rect 553822 588338 587262 588574
rect 587498 588338 587582 588574
rect 587818 588338 592650 588574
rect -8726 588306 592650 588338
rect -8726 585174 592650 585206
rect -8726 584938 -2934 585174
rect -2698 584938 -2614 585174
rect -2378 584938 5546 585174
rect 5782 584938 5866 585174
rect 6102 584938 39546 585174
rect 39782 584938 39866 585174
rect 40102 584938 73546 585174
rect 73782 584938 73866 585174
rect 74102 584938 107546 585174
rect 107782 584938 107866 585174
rect 108102 584938 141546 585174
rect 141782 584938 141866 585174
rect 142102 584938 175546 585174
rect 175782 584938 175866 585174
rect 176102 584938 209546 585174
rect 209782 584938 209866 585174
rect 210102 584938 243546 585174
rect 243782 584938 243866 585174
rect 244102 584938 277546 585174
rect 277782 584938 277866 585174
rect 278102 584938 311546 585174
rect 311782 584938 311866 585174
rect 312102 584938 345546 585174
rect 345782 584938 345866 585174
rect 346102 584938 379546 585174
rect 379782 584938 379866 585174
rect 380102 584938 413546 585174
rect 413782 584938 413866 585174
rect 414102 584938 447546 585174
rect 447782 584938 447866 585174
rect 448102 584938 481546 585174
rect 481782 584938 481866 585174
rect 482102 584938 515546 585174
rect 515782 584938 515866 585174
rect 516102 584938 549546 585174
rect 549782 584938 549866 585174
rect 550102 584938 586302 585174
rect 586538 584938 586622 585174
rect 586858 584938 592650 585174
rect -8726 584854 592650 584938
rect -8726 584618 -2934 584854
rect -2698 584618 -2614 584854
rect -2378 584618 5546 584854
rect 5782 584618 5866 584854
rect 6102 584618 39546 584854
rect 39782 584618 39866 584854
rect 40102 584618 73546 584854
rect 73782 584618 73866 584854
rect 74102 584618 107546 584854
rect 107782 584618 107866 584854
rect 108102 584618 141546 584854
rect 141782 584618 141866 584854
rect 142102 584618 175546 584854
rect 175782 584618 175866 584854
rect 176102 584618 209546 584854
rect 209782 584618 209866 584854
rect 210102 584618 243546 584854
rect 243782 584618 243866 584854
rect 244102 584618 277546 584854
rect 277782 584618 277866 584854
rect 278102 584618 311546 584854
rect 311782 584618 311866 584854
rect 312102 584618 345546 584854
rect 345782 584618 345866 584854
rect 346102 584618 379546 584854
rect 379782 584618 379866 584854
rect 380102 584618 413546 584854
rect 413782 584618 413866 584854
rect 414102 584618 447546 584854
rect 447782 584618 447866 584854
rect 448102 584618 481546 584854
rect 481782 584618 481866 584854
rect 482102 584618 515546 584854
rect 515782 584618 515866 584854
rect 516102 584618 549546 584854
rect 549782 584618 549866 584854
rect 550102 584618 586302 584854
rect 586538 584618 586622 584854
rect 586858 584618 592650 584854
rect -8726 584586 592650 584618
rect -8726 581454 592650 581486
rect -8726 581218 -1974 581454
rect -1738 581218 -1654 581454
rect -1418 581218 1826 581454
rect 2062 581218 2146 581454
rect 2382 581218 35826 581454
rect 36062 581218 36146 581454
rect 36382 581218 69826 581454
rect 70062 581218 70146 581454
rect 70382 581218 103826 581454
rect 104062 581218 104146 581454
rect 104382 581218 137826 581454
rect 138062 581218 138146 581454
rect 138382 581218 171826 581454
rect 172062 581218 172146 581454
rect 172382 581218 205826 581454
rect 206062 581218 206146 581454
rect 206382 581218 239826 581454
rect 240062 581218 240146 581454
rect 240382 581218 273826 581454
rect 274062 581218 274146 581454
rect 274382 581218 307826 581454
rect 308062 581218 308146 581454
rect 308382 581218 341826 581454
rect 342062 581218 342146 581454
rect 342382 581218 375826 581454
rect 376062 581218 376146 581454
rect 376382 581218 409826 581454
rect 410062 581218 410146 581454
rect 410382 581218 443826 581454
rect 444062 581218 444146 581454
rect 444382 581218 477826 581454
rect 478062 581218 478146 581454
rect 478382 581218 511826 581454
rect 512062 581218 512146 581454
rect 512382 581218 545826 581454
rect 546062 581218 546146 581454
rect 546382 581218 579826 581454
rect 580062 581218 580146 581454
rect 580382 581218 585342 581454
rect 585578 581218 585662 581454
rect 585898 581218 592650 581454
rect -8726 581134 592650 581218
rect -8726 580898 -1974 581134
rect -1738 580898 -1654 581134
rect -1418 580898 1826 581134
rect 2062 580898 2146 581134
rect 2382 580898 35826 581134
rect 36062 580898 36146 581134
rect 36382 580898 69826 581134
rect 70062 580898 70146 581134
rect 70382 580898 103826 581134
rect 104062 580898 104146 581134
rect 104382 580898 137826 581134
rect 138062 580898 138146 581134
rect 138382 580898 171826 581134
rect 172062 580898 172146 581134
rect 172382 580898 205826 581134
rect 206062 580898 206146 581134
rect 206382 580898 239826 581134
rect 240062 580898 240146 581134
rect 240382 580898 273826 581134
rect 274062 580898 274146 581134
rect 274382 580898 307826 581134
rect 308062 580898 308146 581134
rect 308382 580898 341826 581134
rect 342062 580898 342146 581134
rect 342382 580898 375826 581134
rect 376062 580898 376146 581134
rect 376382 580898 409826 581134
rect 410062 580898 410146 581134
rect 410382 580898 443826 581134
rect 444062 580898 444146 581134
rect 444382 580898 477826 581134
rect 478062 580898 478146 581134
rect 478382 580898 511826 581134
rect 512062 580898 512146 581134
rect 512382 580898 545826 581134
rect 546062 580898 546146 581134
rect 546382 580898 579826 581134
rect 580062 580898 580146 581134
rect 580382 580898 585342 581134
rect 585578 580898 585662 581134
rect 585898 580898 592650 581134
rect -8726 580866 592650 580898
rect -8726 573494 592650 573526
rect -8726 573258 -8694 573494
rect -8458 573258 -8374 573494
rect -8138 573258 27866 573494
rect 28102 573258 28186 573494
rect 28422 573258 61866 573494
rect 62102 573258 62186 573494
rect 62422 573258 95866 573494
rect 96102 573258 96186 573494
rect 96422 573258 129866 573494
rect 130102 573258 130186 573494
rect 130422 573258 163866 573494
rect 164102 573258 164186 573494
rect 164422 573258 197866 573494
rect 198102 573258 198186 573494
rect 198422 573258 231866 573494
rect 232102 573258 232186 573494
rect 232422 573258 265866 573494
rect 266102 573258 266186 573494
rect 266422 573258 299866 573494
rect 300102 573258 300186 573494
rect 300422 573258 333866 573494
rect 334102 573258 334186 573494
rect 334422 573258 367866 573494
rect 368102 573258 368186 573494
rect 368422 573258 401866 573494
rect 402102 573258 402186 573494
rect 402422 573258 435866 573494
rect 436102 573258 436186 573494
rect 436422 573258 469866 573494
rect 470102 573258 470186 573494
rect 470422 573258 503866 573494
rect 504102 573258 504186 573494
rect 504422 573258 537866 573494
rect 538102 573258 538186 573494
rect 538422 573258 571866 573494
rect 572102 573258 572186 573494
rect 572422 573258 592062 573494
rect 592298 573258 592382 573494
rect 592618 573258 592650 573494
rect -8726 573174 592650 573258
rect -8726 572938 -8694 573174
rect -8458 572938 -8374 573174
rect -8138 572938 27866 573174
rect 28102 572938 28186 573174
rect 28422 572938 61866 573174
rect 62102 572938 62186 573174
rect 62422 572938 95866 573174
rect 96102 572938 96186 573174
rect 96422 572938 129866 573174
rect 130102 572938 130186 573174
rect 130422 572938 163866 573174
rect 164102 572938 164186 573174
rect 164422 572938 197866 573174
rect 198102 572938 198186 573174
rect 198422 572938 231866 573174
rect 232102 572938 232186 573174
rect 232422 572938 265866 573174
rect 266102 572938 266186 573174
rect 266422 572938 299866 573174
rect 300102 572938 300186 573174
rect 300422 572938 333866 573174
rect 334102 572938 334186 573174
rect 334422 572938 367866 573174
rect 368102 572938 368186 573174
rect 368422 572938 401866 573174
rect 402102 572938 402186 573174
rect 402422 572938 435866 573174
rect 436102 572938 436186 573174
rect 436422 572938 469866 573174
rect 470102 572938 470186 573174
rect 470422 572938 503866 573174
rect 504102 572938 504186 573174
rect 504422 572938 537866 573174
rect 538102 572938 538186 573174
rect 538422 572938 571866 573174
rect 572102 572938 572186 573174
rect 572422 572938 592062 573174
rect 592298 572938 592382 573174
rect 592618 572938 592650 573174
rect -8726 572906 592650 572938
rect -8726 569774 592650 569806
rect -8726 569538 -7734 569774
rect -7498 569538 -7414 569774
rect -7178 569538 24146 569774
rect 24382 569538 24466 569774
rect 24702 569538 58146 569774
rect 58382 569538 58466 569774
rect 58702 569538 92146 569774
rect 92382 569538 92466 569774
rect 92702 569538 126146 569774
rect 126382 569538 126466 569774
rect 126702 569538 160146 569774
rect 160382 569538 160466 569774
rect 160702 569538 194146 569774
rect 194382 569538 194466 569774
rect 194702 569538 228146 569774
rect 228382 569538 228466 569774
rect 228702 569538 262146 569774
rect 262382 569538 262466 569774
rect 262702 569538 296146 569774
rect 296382 569538 296466 569774
rect 296702 569538 330146 569774
rect 330382 569538 330466 569774
rect 330702 569538 364146 569774
rect 364382 569538 364466 569774
rect 364702 569538 398146 569774
rect 398382 569538 398466 569774
rect 398702 569538 432146 569774
rect 432382 569538 432466 569774
rect 432702 569538 466146 569774
rect 466382 569538 466466 569774
rect 466702 569538 500146 569774
rect 500382 569538 500466 569774
rect 500702 569538 534146 569774
rect 534382 569538 534466 569774
rect 534702 569538 568146 569774
rect 568382 569538 568466 569774
rect 568702 569538 591102 569774
rect 591338 569538 591422 569774
rect 591658 569538 592650 569774
rect -8726 569454 592650 569538
rect -8726 569218 -7734 569454
rect -7498 569218 -7414 569454
rect -7178 569218 24146 569454
rect 24382 569218 24466 569454
rect 24702 569218 58146 569454
rect 58382 569218 58466 569454
rect 58702 569218 92146 569454
rect 92382 569218 92466 569454
rect 92702 569218 126146 569454
rect 126382 569218 126466 569454
rect 126702 569218 160146 569454
rect 160382 569218 160466 569454
rect 160702 569218 194146 569454
rect 194382 569218 194466 569454
rect 194702 569218 228146 569454
rect 228382 569218 228466 569454
rect 228702 569218 262146 569454
rect 262382 569218 262466 569454
rect 262702 569218 296146 569454
rect 296382 569218 296466 569454
rect 296702 569218 330146 569454
rect 330382 569218 330466 569454
rect 330702 569218 364146 569454
rect 364382 569218 364466 569454
rect 364702 569218 398146 569454
rect 398382 569218 398466 569454
rect 398702 569218 432146 569454
rect 432382 569218 432466 569454
rect 432702 569218 466146 569454
rect 466382 569218 466466 569454
rect 466702 569218 500146 569454
rect 500382 569218 500466 569454
rect 500702 569218 534146 569454
rect 534382 569218 534466 569454
rect 534702 569218 568146 569454
rect 568382 569218 568466 569454
rect 568702 569218 591102 569454
rect 591338 569218 591422 569454
rect 591658 569218 592650 569454
rect -8726 569186 592650 569218
rect -8726 566054 592650 566086
rect -8726 565818 -6774 566054
rect -6538 565818 -6454 566054
rect -6218 565818 20426 566054
rect 20662 565818 20746 566054
rect 20982 565818 54426 566054
rect 54662 565818 54746 566054
rect 54982 565818 88426 566054
rect 88662 565818 88746 566054
rect 88982 565818 122426 566054
rect 122662 565818 122746 566054
rect 122982 565818 156426 566054
rect 156662 565818 156746 566054
rect 156982 565818 190426 566054
rect 190662 565818 190746 566054
rect 190982 565818 224426 566054
rect 224662 565818 224746 566054
rect 224982 565818 258426 566054
rect 258662 565818 258746 566054
rect 258982 565818 292426 566054
rect 292662 565818 292746 566054
rect 292982 565818 326426 566054
rect 326662 565818 326746 566054
rect 326982 565818 360426 566054
rect 360662 565818 360746 566054
rect 360982 565818 394426 566054
rect 394662 565818 394746 566054
rect 394982 565818 428426 566054
rect 428662 565818 428746 566054
rect 428982 565818 462426 566054
rect 462662 565818 462746 566054
rect 462982 565818 496426 566054
rect 496662 565818 496746 566054
rect 496982 565818 530426 566054
rect 530662 565818 530746 566054
rect 530982 565818 564426 566054
rect 564662 565818 564746 566054
rect 564982 565818 590142 566054
rect 590378 565818 590462 566054
rect 590698 565818 592650 566054
rect -8726 565734 592650 565818
rect -8726 565498 -6774 565734
rect -6538 565498 -6454 565734
rect -6218 565498 20426 565734
rect 20662 565498 20746 565734
rect 20982 565498 54426 565734
rect 54662 565498 54746 565734
rect 54982 565498 88426 565734
rect 88662 565498 88746 565734
rect 88982 565498 122426 565734
rect 122662 565498 122746 565734
rect 122982 565498 156426 565734
rect 156662 565498 156746 565734
rect 156982 565498 190426 565734
rect 190662 565498 190746 565734
rect 190982 565498 224426 565734
rect 224662 565498 224746 565734
rect 224982 565498 258426 565734
rect 258662 565498 258746 565734
rect 258982 565498 292426 565734
rect 292662 565498 292746 565734
rect 292982 565498 326426 565734
rect 326662 565498 326746 565734
rect 326982 565498 360426 565734
rect 360662 565498 360746 565734
rect 360982 565498 394426 565734
rect 394662 565498 394746 565734
rect 394982 565498 428426 565734
rect 428662 565498 428746 565734
rect 428982 565498 462426 565734
rect 462662 565498 462746 565734
rect 462982 565498 496426 565734
rect 496662 565498 496746 565734
rect 496982 565498 530426 565734
rect 530662 565498 530746 565734
rect 530982 565498 564426 565734
rect 564662 565498 564746 565734
rect 564982 565498 590142 565734
rect 590378 565498 590462 565734
rect 590698 565498 592650 565734
rect -8726 565466 592650 565498
rect -8726 562334 592650 562366
rect -8726 562098 -5814 562334
rect -5578 562098 -5494 562334
rect -5258 562098 16706 562334
rect 16942 562098 17026 562334
rect 17262 562098 50706 562334
rect 50942 562098 51026 562334
rect 51262 562098 84706 562334
rect 84942 562098 85026 562334
rect 85262 562098 118706 562334
rect 118942 562098 119026 562334
rect 119262 562098 152706 562334
rect 152942 562098 153026 562334
rect 153262 562098 186706 562334
rect 186942 562098 187026 562334
rect 187262 562098 220706 562334
rect 220942 562098 221026 562334
rect 221262 562098 254706 562334
rect 254942 562098 255026 562334
rect 255262 562098 288706 562334
rect 288942 562098 289026 562334
rect 289262 562098 322706 562334
rect 322942 562098 323026 562334
rect 323262 562098 356706 562334
rect 356942 562098 357026 562334
rect 357262 562098 390706 562334
rect 390942 562098 391026 562334
rect 391262 562098 424706 562334
rect 424942 562098 425026 562334
rect 425262 562098 458706 562334
rect 458942 562098 459026 562334
rect 459262 562098 492706 562334
rect 492942 562098 493026 562334
rect 493262 562098 526706 562334
rect 526942 562098 527026 562334
rect 527262 562098 560706 562334
rect 560942 562098 561026 562334
rect 561262 562098 589182 562334
rect 589418 562098 589502 562334
rect 589738 562098 592650 562334
rect -8726 562014 592650 562098
rect -8726 561778 -5814 562014
rect -5578 561778 -5494 562014
rect -5258 561778 16706 562014
rect 16942 561778 17026 562014
rect 17262 561778 50706 562014
rect 50942 561778 51026 562014
rect 51262 561778 84706 562014
rect 84942 561778 85026 562014
rect 85262 561778 118706 562014
rect 118942 561778 119026 562014
rect 119262 561778 152706 562014
rect 152942 561778 153026 562014
rect 153262 561778 186706 562014
rect 186942 561778 187026 562014
rect 187262 561778 220706 562014
rect 220942 561778 221026 562014
rect 221262 561778 254706 562014
rect 254942 561778 255026 562014
rect 255262 561778 288706 562014
rect 288942 561778 289026 562014
rect 289262 561778 322706 562014
rect 322942 561778 323026 562014
rect 323262 561778 356706 562014
rect 356942 561778 357026 562014
rect 357262 561778 390706 562014
rect 390942 561778 391026 562014
rect 391262 561778 424706 562014
rect 424942 561778 425026 562014
rect 425262 561778 458706 562014
rect 458942 561778 459026 562014
rect 459262 561778 492706 562014
rect 492942 561778 493026 562014
rect 493262 561778 526706 562014
rect 526942 561778 527026 562014
rect 527262 561778 560706 562014
rect 560942 561778 561026 562014
rect 561262 561778 589182 562014
rect 589418 561778 589502 562014
rect 589738 561778 592650 562014
rect -8726 561746 592650 561778
rect -8726 558614 592650 558646
rect -8726 558378 -4854 558614
rect -4618 558378 -4534 558614
rect -4298 558378 12986 558614
rect 13222 558378 13306 558614
rect 13542 558378 46986 558614
rect 47222 558378 47306 558614
rect 47542 558378 80986 558614
rect 81222 558378 81306 558614
rect 81542 558378 114986 558614
rect 115222 558378 115306 558614
rect 115542 558378 148986 558614
rect 149222 558378 149306 558614
rect 149542 558378 182986 558614
rect 183222 558378 183306 558614
rect 183542 558378 216986 558614
rect 217222 558378 217306 558614
rect 217542 558378 250986 558614
rect 251222 558378 251306 558614
rect 251542 558378 284986 558614
rect 285222 558378 285306 558614
rect 285542 558378 318986 558614
rect 319222 558378 319306 558614
rect 319542 558378 352986 558614
rect 353222 558378 353306 558614
rect 353542 558378 386986 558614
rect 387222 558378 387306 558614
rect 387542 558378 420986 558614
rect 421222 558378 421306 558614
rect 421542 558378 454986 558614
rect 455222 558378 455306 558614
rect 455542 558378 488986 558614
rect 489222 558378 489306 558614
rect 489542 558378 522986 558614
rect 523222 558378 523306 558614
rect 523542 558378 556986 558614
rect 557222 558378 557306 558614
rect 557542 558378 588222 558614
rect 588458 558378 588542 558614
rect 588778 558378 592650 558614
rect -8726 558294 592650 558378
rect -8726 558058 -4854 558294
rect -4618 558058 -4534 558294
rect -4298 558058 12986 558294
rect 13222 558058 13306 558294
rect 13542 558058 46986 558294
rect 47222 558058 47306 558294
rect 47542 558058 80986 558294
rect 81222 558058 81306 558294
rect 81542 558058 114986 558294
rect 115222 558058 115306 558294
rect 115542 558058 148986 558294
rect 149222 558058 149306 558294
rect 149542 558058 182986 558294
rect 183222 558058 183306 558294
rect 183542 558058 216986 558294
rect 217222 558058 217306 558294
rect 217542 558058 250986 558294
rect 251222 558058 251306 558294
rect 251542 558058 284986 558294
rect 285222 558058 285306 558294
rect 285542 558058 318986 558294
rect 319222 558058 319306 558294
rect 319542 558058 352986 558294
rect 353222 558058 353306 558294
rect 353542 558058 386986 558294
rect 387222 558058 387306 558294
rect 387542 558058 420986 558294
rect 421222 558058 421306 558294
rect 421542 558058 454986 558294
rect 455222 558058 455306 558294
rect 455542 558058 488986 558294
rect 489222 558058 489306 558294
rect 489542 558058 522986 558294
rect 523222 558058 523306 558294
rect 523542 558058 556986 558294
rect 557222 558058 557306 558294
rect 557542 558058 588222 558294
rect 588458 558058 588542 558294
rect 588778 558058 592650 558294
rect -8726 558026 592650 558058
rect -8726 554894 592650 554926
rect -8726 554658 -3894 554894
rect -3658 554658 -3574 554894
rect -3338 554658 9266 554894
rect 9502 554658 9586 554894
rect 9822 554658 43266 554894
rect 43502 554658 43586 554894
rect 43822 554658 77266 554894
rect 77502 554658 77586 554894
rect 77822 554658 111266 554894
rect 111502 554658 111586 554894
rect 111822 554658 145266 554894
rect 145502 554658 145586 554894
rect 145822 554658 179266 554894
rect 179502 554658 179586 554894
rect 179822 554658 213266 554894
rect 213502 554658 213586 554894
rect 213822 554658 247266 554894
rect 247502 554658 247586 554894
rect 247822 554658 281266 554894
rect 281502 554658 281586 554894
rect 281822 554658 315266 554894
rect 315502 554658 315586 554894
rect 315822 554658 349266 554894
rect 349502 554658 349586 554894
rect 349822 554658 383266 554894
rect 383502 554658 383586 554894
rect 383822 554658 417266 554894
rect 417502 554658 417586 554894
rect 417822 554658 451266 554894
rect 451502 554658 451586 554894
rect 451822 554658 485266 554894
rect 485502 554658 485586 554894
rect 485822 554658 519266 554894
rect 519502 554658 519586 554894
rect 519822 554658 553266 554894
rect 553502 554658 553586 554894
rect 553822 554658 587262 554894
rect 587498 554658 587582 554894
rect 587818 554658 592650 554894
rect -8726 554574 592650 554658
rect -8726 554338 -3894 554574
rect -3658 554338 -3574 554574
rect -3338 554338 9266 554574
rect 9502 554338 9586 554574
rect 9822 554338 43266 554574
rect 43502 554338 43586 554574
rect 43822 554338 77266 554574
rect 77502 554338 77586 554574
rect 77822 554338 111266 554574
rect 111502 554338 111586 554574
rect 111822 554338 145266 554574
rect 145502 554338 145586 554574
rect 145822 554338 179266 554574
rect 179502 554338 179586 554574
rect 179822 554338 213266 554574
rect 213502 554338 213586 554574
rect 213822 554338 247266 554574
rect 247502 554338 247586 554574
rect 247822 554338 281266 554574
rect 281502 554338 281586 554574
rect 281822 554338 315266 554574
rect 315502 554338 315586 554574
rect 315822 554338 349266 554574
rect 349502 554338 349586 554574
rect 349822 554338 383266 554574
rect 383502 554338 383586 554574
rect 383822 554338 417266 554574
rect 417502 554338 417586 554574
rect 417822 554338 451266 554574
rect 451502 554338 451586 554574
rect 451822 554338 485266 554574
rect 485502 554338 485586 554574
rect 485822 554338 519266 554574
rect 519502 554338 519586 554574
rect 519822 554338 553266 554574
rect 553502 554338 553586 554574
rect 553822 554338 587262 554574
rect 587498 554338 587582 554574
rect 587818 554338 592650 554574
rect -8726 554306 592650 554338
rect -8726 551174 592650 551206
rect -8726 550938 -2934 551174
rect -2698 550938 -2614 551174
rect -2378 550938 5546 551174
rect 5782 550938 5866 551174
rect 6102 550938 39546 551174
rect 39782 550938 39866 551174
rect 40102 550938 73546 551174
rect 73782 550938 73866 551174
rect 74102 550938 107546 551174
rect 107782 550938 107866 551174
rect 108102 550938 141546 551174
rect 141782 550938 141866 551174
rect 142102 550938 175546 551174
rect 175782 550938 175866 551174
rect 176102 550938 209546 551174
rect 209782 550938 209866 551174
rect 210102 550938 243546 551174
rect 243782 550938 243866 551174
rect 244102 550938 277546 551174
rect 277782 550938 277866 551174
rect 278102 550938 311546 551174
rect 311782 550938 311866 551174
rect 312102 550938 345546 551174
rect 345782 550938 345866 551174
rect 346102 550938 379546 551174
rect 379782 550938 379866 551174
rect 380102 550938 413546 551174
rect 413782 550938 413866 551174
rect 414102 550938 447546 551174
rect 447782 550938 447866 551174
rect 448102 550938 481546 551174
rect 481782 550938 481866 551174
rect 482102 550938 515546 551174
rect 515782 550938 515866 551174
rect 516102 550938 549546 551174
rect 549782 550938 549866 551174
rect 550102 550938 586302 551174
rect 586538 550938 586622 551174
rect 586858 550938 592650 551174
rect -8726 550854 592650 550938
rect -8726 550618 -2934 550854
rect -2698 550618 -2614 550854
rect -2378 550618 5546 550854
rect 5782 550618 5866 550854
rect 6102 550618 39546 550854
rect 39782 550618 39866 550854
rect 40102 550618 73546 550854
rect 73782 550618 73866 550854
rect 74102 550618 107546 550854
rect 107782 550618 107866 550854
rect 108102 550618 141546 550854
rect 141782 550618 141866 550854
rect 142102 550618 175546 550854
rect 175782 550618 175866 550854
rect 176102 550618 209546 550854
rect 209782 550618 209866 550854
rect 210102 550618 243546 550854
rect 243782 550618 243866 550854
rect 244102 550618 277546 550854
rect 277782 550618 277866 550854
rect 278102 550618 311546 550854
rect 311782 550618 311866 550854
rect 312102 550618 345546 550854
rect 345782 550618 345866 550854
rect 346102 550618 379546 550854
rect 379782 550618 379866 550854
rect 380102 550618 413546 550854
rect 413782 550618 413866 550854
rect 414102 550618 447546 550854
rect 447782 550618 447866 550854
rect 448102 550618 481546 550854
rect 481782 550618 481866 550854
rect 482102 550618 515546 550854
rect 515782 550618 515866 550854
rect 516102 550618 549546 550854
rect 549782 550618 549866 550854
rect 550102 550618 586302 550854
rect 586538 550618 586622 550854
rect 586858 550618 592650 550854
rect -8726 550586 592650 550618
rect -8726 547454 592650 547486
rect -8726 547218 -1974 547454
rect -1738 547218 -1654 547454
rect -1418 547218 1826 547454
rect 2062 547218 2146 547454
rect 2382 547218 35826 547454
rect 36062 547218 36146 547454
rect 36382 547218 69826 547454
rect 70062 547218 70146 547454
rect 70382 547218 103826 547454
rect 104062 547218 104146 547454
rect 104382 547218 137826 547454
rect 138062 547218 138146 547454
rect 138382 547218 171826 547454
rect 172062 547218 172146 547454
rect 172382 547218 205826 547454
rect 206062 547218 206146 547454
rect 206382 547218 239826 547454
rect 240062 547218 240146 547454
rect 240382 547218 273826 547454
rect 274062 547218 274146 547454
rect 274382 547218 307826 547454
rect 308062 547218 308146 547454
rect 308382 547218 341826 547454
rect 342062 547218 342146 547454
rect 342382 547218 375826 547454
rect 376062 547218 376146 547454
rect 376382 547218 409826 547454
rect 410062 547218 410146 547454
rect 410382 547218 443826 547454
rect 444062 547218 444146 547454
rect 444382 547218 477826 547454
rect 478062 547218 478146 547454
rect 478382 547218 511826 547454
rect 512062 547218 512146 547454
rect 512382 547218 545826 547454
rect 546062 547218 546146 547454
rect 546382 547218 579826 547454
rect 580062 547218 580146 547454
rect 580382 547218 585342 547454
rect 585578 547218 585662 547454
rect 585898 547218 592650 547454
rect -8726 547134 592650 547218
rect -8726 546898 -1974 547134
rect -1738 546898 -1654 547134
rect -1418 546898 1826 547134
rect 2062 546898 2146 547134
rect 2382 546898 35826 547134
rect 36062 546898 36146 547134
rect 36382 546898 69826 547134
rect 70062 546898 70146 547134
rect 70382 546898 103826 547134
rect 104062 546898 104146 547134
rect 104382 546898 137826 547134
rect 138062 546898 138146 547134
rect 138382 546898 171826 547134
rect 172062 546898 172146 547134
rect 172382 546898 205826 547134
rect 206062 546898 206146 547134
rect 206382 546898 239826 547134
rect 240062 546898 240146 547134
rect 240382 546898 273826 547134
rect 274062 546898 274146 547134
rect 274382 546898 307826 547134
rect 308062 546898 308146 547134
rect 308382 546898 341826 547134
rect 342062 546898 342146 547134
rect 342382 546898 375826 547134
rect 376062 546898 376146 547134
rect 376382 546898 409826 547134
rect 410062 546898 410146 547134
rect 410382 546898 443826 547134
rect 444062 546898 444146 547134
rect 444382 546898 477826 547134
rect 478062 546898 478146 547134
rect 478382 546898 511826 547134
rect 512062 546898 512146 547134
rect 512382 546898 545826 547134
rect 546062 546898 546146 547134
rect 546382 546898 579826 547134
rect 580062 546898 580146 547134
rect 580382 546898 585342 547134
rect 585578 546898 585662 547134
rect 585898 546898 592650 547134
rect -8726 546866 592650 546898
rect -8726 539494 592650 539526
rect -8726 539258 -8694 539494
rect -8458 539258 -8374 539494
rect -8138 539258 27866 539494
rect 28102 539258 28186 539494
rect 28422 539258 61866 539494
rect 62102 539258 62186 539494
rect 62422 539258 95866 539494
rect 96102 539258 96186 539494
rect 96422 539258 129866 539494
rect 130102 539258 130186 539494
rect 130422 539258 163866 539494
rect 164102 539258 164186 539494
rect 164422 539258 197866 539494
rect 198102 539258 198186 539494
rect 198422 539258 231866 539494
rect 232102 539258 232186 539494
rect 232422 539258 265866 539494
rect 266102 539258 266186 539494
rect 266422 539258 299866 539494
rect 300102 539258 300186 539494
rect 300422 539258 333866 539494
rect 334102 539258 334186 539494
rect 334422 539258 367866 539494
rect 368102 539258 368186 539494
rect 368422 539258 401866 539494
rect 402102 539258 402186 539494
rect 402422 539258 435866 539494
rect 436102 539258 436186 539494
rect 436422 539258 469866 539494
rect 470102 539258 470186 539494
rect 470422 539258 503866 539494
rect 504102 539258 504186 539494
rect 504422 539258 537866 539494
rect 538102 539258 538186 539494
rect 538422 539258 571866 539494
rect 572102 539258 572186 539494
rect 572422 539258 592062 539494
rect 592298 539258 592382 539494
rect 592618 539258 592650 539494
rect -8726 539174 592650 539258
rect -8726 538938 -8694 539174
rect -8458 538938 -8374 539174
rect -8138 538938 27866 539174
rect 28102 538938 28186 539174
rect 28422 538938 61866 539174
rect 62102 538938 62186 539174
rect 62422 538938 95866 539174
rect 96102 538938 96186 539174
rect 96422 538938 129866 539174
rect 130102 538938 130186 539174
rect 130422 538938 163866 539174
rect 164102 538938 164186 539174
rect 164422 538938 197866 539174
rect 198102 538938 198186 539174
rect 198422 538938 231866 539174
rect 232102 538938 232186 539174
rect 232422 538938 265866 539174
rect 266102 538938 266186 539174
rect 266422 538938 299866 539174
rect 300102 538938 300186 539174
rect 300422 538938 333866 539174
rect 334102 538938 334186 539174
rect 334422 538938 367866 539174
rect 368102 538938 368186 539174
rect 368422 538938 401866 539174
rect 402102 538938 402186 539174
rect 402422 538938 435866 539174
rect 436102 538938 436186 539174
rect 436422 538938 469866 539174
rect 470102 538938 470186 539174
rect 470422 538938 503866 539174
rect 504102 538938 504186 539174
rect 504422 538938 537866 539174
rect 538102 538938 538186 539174
rect 538422 538938 571866 539174
rect 572102 538938 572186 539174
rect 572422 538938 592062 539174
rect 592298 538938 592382 539174
rect 592618 538938 592650 539174
rect -8726 538906 592650 538938
rect -8726 535774 592650 535806
rect -8726 535538 -7734 535774
rect -7498 535538 -7414 535774
rect -7178 535538 24146 535774
rect 24382 535538 24466 535774
rect 24702 535538 58146 535774
rect 58382 535538 58466 535774
rect 58702 535538 92146 535774
rect 92382 535538 92466 535774
rect 92702 535538 126146 535774
rect 126382 535538 126466 535774
rect 126702 535538 160146 535774
rect 160382 535538 160466 535774
rect 160702 535538 194146 535774
rect 194382 535538 194466 535774
rect 194702 535538 228146 535774
rect 228382 535538 228466 535774
rect 228702 535538 262146 535774
rect 262382 535538 262466 535774
rect 262702 535538 296146 535774
rect 296382 535538 296466 535774
rect 296702 535538 330146 535774
rect 330382 535538 330466 535774
rect 330702 535538 364146 535774
rect 364382 535538 364466 535774
rect 364702 535538 398146 535774
rect 398382 535538 398466 535774
rect 398702 535538 432146 535774
rect 432382 535538 432466 535774
rect 432702 535538 466146 535774
rect 466382 535538 466466 535774
rect 466702 535538 500146 535774
rect 500382 535538 500466 535774
rect 500702 535538 534146 535774
rect 534382 535538 534466 535774
rect 534702 535538 568146 535774
rect 568382 535538 568466 535774
rect 568702 535538 591102 535774
rect 591338 535538 591422 535774
rect 591658 535538 592650 535774
rect -8726 535454 592650 535538
rect -8726 535218 -7734 535454
rect -7498 535218 -7414 535454
rect -7178 535218 24146 535454
rect 24382 535218 24466 535454
rect 24702 535218 58146 535454
rect 58382 535218 58466 535454
rect 58702 535218 92146 535454
rect 92382 535218 92466 535454
rect 92702 535218 126146 535454
rect 126382 535218 126466 535454
rect 126702 535218 160146 535454
rect 160382 535218 160466 535454
rect 160702 535218 194146 535454
rect 194382 535218 194466 535454
rect 194702 535218 228146 535454
rect 228382 535218 228466 535454
rect 228702 535218 262146 535454
rect 262382 535218 262466 535454
rect 262702 535218 296146 535454
rect 296382 535218 296466 535454
rect 296702 535218 330146 535454
rect 330382 535218 330466 535454
rect 330702 535218 364146 535454
rect 364382 535218 364466 535454
rect 364702 535218 398146 535454
rect 398382 535218 398466 535454
rect 398702 535218 432146 535454
rect 432382 535218 432466 535454
rect 432702 535218 466146 535454
rect 466382 535218 466466 535454
rect 466702 535218 500146 535454
rect 500382 535218 500466 535454
rect 500702 535218 534146 535454
rect 534382 535218 534466 535454
rect 534702 535218 568146 535454
rect 568382 535218 568466 535454
rect 568702 535218 591102 535454
rect 591338 535218 591422 535454
rect 591658 535218 592650 535454
rect -8726 535186 592650 535218
rect -8726 532054 592650 532086
rect -8726 531818 -6774 532054
rect -6538 531818 -6454 532054
rect -6218 531818 20426 532054
rect 20662 531818 20746 532054
rect 20982 531818 54426 532054
rect 54662 531818 54746 532054
rect 54982 531818 88426 532054
rect 88662 531818 88746 532054
rect 88982 531818 122426 532054
rect 122662 531818 122746 532054
rect 122982 531818 156426 532054
rect 156662 531818 156746 532054
rect 156982 531818 190426 532054
rect 190662 531818 190746 532054
rect 190982 531818 224426 532054
rect 224662 531818 224746 532054
rect 224982 531818 258426 532054
rect 258662 531818 258746 532054
rect 258982 531818 292426 532054
rect 292662 531818 292746 532054
rect 292982 531818 326426 532054
rect 326662 531818 326746 532054
rect 326982 531818 360426 532054
rect 360662 531818 360746 532054
rect 360982 531818 394426 532054
rect 394662 531818 394746 532054
rect 394982 531818 428426 532054
rect 428662 531818 428746 532054
rect 428982 531818 462426 532054
rect 462662 531818 462746 532054
rect 462982 531818 496426 532054
rect 496662 531818 496746 532054
rect 496982 531818 530426 532054
rect 530662 531818 530746 532054
rect 530982 531818 564426 532054
rect 564662 531818 564746 532054
rect 564982 531818 590142 532054
rect 590378 531818 590462 532054
rect 590698 531818 592650 532054
rect -8726 531734 592650 531818
rect -8726 531498 -6774 531734
rect -6538 531498 -6454 531734
rect -6218 531498 20426 531734
rect 20662 531498 20746 531734
rect 20982 531498 54426 531734
rect 54662 531498 54746 531734
rect 54982 531498 88426 531734
rect 88662 531498 88746 531734
rect 88982 531498 122426 531734
rect 122662 531498 122746 531734
rect 122982 531498 156426 531734
rect 156662 531498 156746 531734
rect 156982 531498 190426 531734
rect 190662 531498 190746 531734
rect 190982 531498 224426 531734
rect 224662 531498 224746 531734
rect 224982 531498 258426 531734
rect 258662 531498 258746 531734
rect 258982 531498 292426 531734
rect 292662 531498 292746 531734
rect 292982 531498 326426 531734
rect 326662 531498 326746 531734
rect 326982 531498 360426 531734
rect 360662 531498 360746 531734
rect 360982 531498 394426 531734
rect 394662 531498 394746 531734
rect 394982 531498 428426 531734
rect 428662 531498 428746 531734
rect 428982 531498 462426 531734
rect 462662 531498 462746 531734
rect 462982 531498 496426 531734
rect 496662 531498 496746 531734
rect 496982 531498 530426 531734
rect 530662 531498 530746 531734
rect 530982 531498 564426 531734
rect 564662 531498 564746 531734
rect 564982 531498 590142 531734
rect 590378 531498 590462 531734
rect 590698 531498 592650 531734
rect -8726 531466 592650 531498
rect -8726 528334 592650 528366
rect -8726 528098 -5814 528334
rect -5578 528098 -5494 528334
rect -5258 528098 16706 528334
rect 16942 528098 17026 528334
rect 17262 528098 50706 528334
rect 50942 528098 51026 528334
rect 51262 528098 84706 528334
rect 84942 528098 85026 528334
rect 85262 528098 118706 528334
rect 118942 528098 119026 528334
rect 119262 528098 152706 528334
rect 152942 528098 153026 528334
rect 153262 528098 186706 528334
rect 186942 528098 187026 528334
rect 187262 528098 220706 528334
rect 220942 528098 221026 528334
rect 221262 528098 254706 528334
rect 254942 528098 255026 528334
rect 255262 528098 288706 528334
rect 288942 528098 289026 528334
rect 289262 528098 322706 528334
rect 322942 528098 323026 528334
rect 323262 528098 356706 528334
rect 356942 528098 357026 528334
rect 357262 528098 390706 528334
rect 390942 528098 391026 528334
rect 391262 528098 424706 528334
rect 424942 528098 425026 528334
rect 425262 528098 458706 528334
rect 458942 528098 459026 528334
rect 459262 528098 492706 528334
rect 492942 528098 493026 528334
rect 493262 528098 526706 528334
rect 526942 528098 527026 528334
rect 527262 528098 560706 528334
rect 560942 528098 561026 528334
rect 561262 528098 589182 528334
rect 589418 528098 589502 528334
rect 589738 528098 592650 528334
rect -8726 528014 592650 528098
rect -8726 527778 -5814 528014
rect -5578 527778 -5494 528014
rect -5258 527778 16706 528014
rect 16942 527778 17026 528014
rect 17262 527778 50706 528014
rect 50942 527778 51026 528014
rect 51262 527778 84706 528014
rect 84942 527778 85026 528014
rect 85262 527778 118706 528014
rect 118942 527778 119026 528014
rect 119262 527778 152706 528014
rect 152942 527778 153026 528014
rect 153262 527778 186706 528014
rect 186942 527778 187026 528014
rect 187262 527778 220706 528014
rect 220942 527778 221026 528014
rect 221262 527778 254706 528014
rect 254942 527778 255026 528014
rect 255262 527778 288706 528014
rect 288942 527778 289026 528014
rect 289262 527778 322706 528014
rect 322942 527778 323026 528014
rect 323262 527778 356706 528014
rect 356942 527778 357026 528014
rect 357262 527778 390706 528014
rect 390942 527778 391026 528014
rect 391262 527778 424706 528014
rect 424942 527778 425026 528014
rect 425262 527778 458706 528014
rect 458942 527778 459026 528014
rect 459262 527778 492706 528014
rect 492942 527778 493026 528014
rect 493262 527778 526706 528014
rect 526942 527778 527026 528014
rect 527262 527778 560706 528014
rect 560942 527778 561026 528014
rect 561262 527778 589182 528014
rect 589418 527778 589502 528014
rect 589738 527778 592650 528014
rect -8726 527746 592650 527778
rect -8726 524614 592650 524646
rect -8726 524378 -4854 524614
rect -4618 524378 -4534 524614
rect -4298 524378 12986 524614
rect 13222 524378 13306 524614
rect 13542 524378 46986 524614
rect 47222 524378 47306 524614
rect 47542 524378 80986 524614
rect 81222 524378 81306 524614
rect 81542 524378 114986 524614
rect 115222 524378 115306 524614
rect 115542 524378 148986 524614
rect 149222 524378 149306 524614
rect 149542 524378 182986 524614
rect 183222 524378 183306 524614
rect 183542 524378 216986 524614
rect 217222 524378 217306 524614
rect 217542 524378 250986 524614
rect 251222 524378 251306 524614
rect 251542 524378 284986 524614
rect 285222 524378 285306 524614
rect 285542 524378 318986 524614
rect 319222 524378 319306 524614
rect 319542 524378 352986 524614
rect 353222 524378 353306 524614
rect 353542 524378 386986 524614
rect 387222 524378 387306 524614
rect 387542 524378 420986 524614
rect 421222 524378 421306 524614
rect 421542 524378 454986 524614
rect 455222 524378 455306 524614
rect 455542 524378 488986 524614
rect 489222 524378 489306 524614
rect 489542 524378 522986 524614
rect 523222 524378 523306 524614
rect 523542 524378 556986 524614
rect 557222 524378 557306 524614
rect 557542 524378 588222 524614
rect 588458 524378 588542 524614
rect 588778 524378 592650 524614
rect -8726 524294 592650 524378
rect -8726 524058 -4854 524294
rect -4618 524058 -4534 524294
rect -4298 524058 12986 524294
rect 13222 524058 13306 524294
rect 13542 524058 46986 524294
rect 47222 524058 47306 524294
rect 47542 524058 80986 524294
rect 81222 524058 81306 524294
rect 81542 524058 114986 524294
rect 115222 524058 115306 524294
rect 115542 524058 148986 524294
rect 149222 524058 149306 524294
rect 149542 524058 182986 524294
rect 183222 524058 183306 524294
rect 183542 524058 216986 524294
rect 217222 524058 217306 524294
rect 217542 524058 250986 524294
rect 251222 524058 251306 524294
rect 251542 524058 284986 524294
rect 285222 524058 285306 524294
rect 285542 524058 318986 524294
rect 319222 524058 319306 524294
rect 319542 524058 352986 524294
rect 353222 524058 353306 524294
rect 353542 524058 386986 524294
rect 387222 524058 387306 524294
rect 387542 524058 420986 524294
rect 421222 524058 421306 524294
rect 421542 524058 454986 524294
rect 455222 524058 455306 524294
rect 455542 524058 488986 524294
rect 489222 524058 489306 524294
rect 489542 524058 522986 524294
rect 523222 524058 523306 524294
rect 523542 524058 556986 524294
rect 557222 524058 557306 524294
rect 557542 524058 588222 524294
rect 588458 524058 588542 524294
rect 588778 524058 592650 524294
rect -8726 524026 592650 524058
rect -8726 520894 592650 520926
rect -8726 520658 -3894 520894
rect -3658 520658 -3574 520894
rect -3338 520658 9266 520894
rect 9502 520658 9586 520894
rect 9822 520658 43266 520894
rect 43502 520658 43586 520894
rect 43822 520658 77266 520894
rect 77502 520658 77586 520894
rect 77822 520658 111266 520894
rect 111502 520658 111586 520894
rect 111822 520658 145266 520894
rect 145502 520658 145586 520894
rect 145822 520658 179266 520894
rect 179502 520658 179586 520894
rect 179822 520658 213266 520894
rect 213502 520658 213586 520894
rect 213822 520658 247266 520894
rect 247502 520658 247586 520894
rect 247822 520658 281266 520894
rect 281502 520658 281586 520894
rect 281822 520658 315266 520894
rect 315502 520658 315586 520894
rect 315822 520658 349266 520894
rect 349502 520658 349586 520894
rect 349822 520658 383266 520894
rect 383502 520658 383586 520894
rect 383822 520658 417266 520894
rect 417502 520658 417586 520894
rect 417822 520658 451266 520894
rect 451502 520658 451586 520894
rect 451822 520658 485266 520894
rect 485502 520658 485586 520894
rect 485822 520658 519266 520894
rect 519502 520658 519586 520894
rect 519822 520658 553266 520894
rect 553502 520658 553586 520894
rect 553822 520658 587262 520894
rect 587498 520658 587582 520894
rect 587818 520658 592650 520894
rect -8726 520574 592650 520658
rect -8726 520338 -3894 520574
rect -3658 520338 -3574 520574
rect -3338 520338 9266 520574
rect 9502 520338 9586 520574
rect 9822 520338 43266 520574
rect 43502 520338 43586 520574
rect 43822 520338 77266 520574
rect 77502 520338 77586 520574
rect 77822 520338 111266 520574
rect 111502 520338 111586 520574
rect 111822 520338 145266 520574
rect 145502 520338 145586 520574
rect 145822 520338 179266 520574
rect 179502 520338 179586 520574
rect 179822 520338 213266 520574
rect 213502 520338 213586 520574
rect 213822 520338 247266 520574
rect 247502 520338 247586 520574
rect 247822 520338 281266 520574
rect 281502 520338 281586 520574
rect 281822 520338 315266 520574
rect 315502 520338 315586 520574
rect 315822 520338 349266 520574
rect 349502 520338 349586 520574
rect 349822 520338 383266 520574
rect 383502 520338 383586 520574
rect 383822 520338 417266 520574
rect 417502 520338 417586 520574
rect 417822 520338 451266 520574
rect 451502 520338 451586 520574
rect 451822 520338 485266 520574
rect 485502 520338 485586 520574
rect 485822 520338 519266 520574
rect 519502 520338 519586 520574
rect 519822 520338 553266 520574
rect 553502 520338 553586 520574
rect 553822 520338 587262 520574
rect 587498 520338 587582 520574
rect 587818 520338 592650 520574
rect -8726 520306 592650 520338
rect -8726 517174 592650 517206
rect -8726 516938 -2934 517174
rect -2698 516938 -2614 517174
rect -2378 516938 5546 517174
rect 5782 516938 5866 517174
rect 6102 516938 39546 517174
rect 39782 516938 39866 517174
rect 40102 516938 73546 517174
rect 73782 516938 73866 517174
rect 74102 516938 107546 517174
rect 107782 516938 107866 517174
rect 108102 516938 141546 517174
rect 141782 516938 141866 517174
rect 142102 516938 175546 517174
rect 175782 516938 175866 517174
rect 176102 516938 209546 517174
rect 209782 516938 209866 517174
rect 210102 516938 243546 517174
rect 243782 516938 243866 517174
rect 244102 516938 277546 517174
rect 277782 516938 277866 517174
rect 278102 516938 311546 517174
rect 311782 516938 311866 517174
rect 312102 516938 345546 517174
rect 345782 516938 345866 517174
rect 346102 516938 379546 517174
rect 379782 516938 379866 517174
rect 380102 516938 413546 517174
rect 413782 516938 413866 517174
rect 414102 516938 447546 517174
rect 447782 516938 447866 517174
rect 448102 516938 481546 517174
rect 481782 516938 481866 517174
rect 482102 516938 515546 517174
rect 515782 516938 515866 517174
rect 516102 516938 549546 517174
rect 549782 516938 549866 517174
rect 550102 516938 586302 517174
rect 586538 516938 586622 517174
rect 586858 516938 592650 517174
rect -8726 516854 592650 516938
rect -8726 516618 -2934 516854
rect -2698 516618 -2614 516854
rect -2378 516618 5546 516854
rect 5782 516618 5866 516854
rect 6102 516618 39546 516854
rect 39782 516618 39866 516854
rect 40102 516618 73546 516854
rect 73782 516618 73866 516854
rect 74102 516618 107546 516854
rect 107782 516618 107866 516854
rect 108102 516618 141546 516854
rect 141782 516618 141866 516854
rect 142102 516618 175546 516854
rect 175782 516618 175866 516854
rect 176102 516618 209546 516854
rect 209782 516618 209866 516854
rect 210102 516618 243546 516854
rect 243782 516618 243866 516854
rect 244102 516618 277546 516854
rect 277782 516618 277866 516854
rect 278102 516618 311546 516854
rect 311782 516618 311866 516854
rect 312102 516618 345546 516854
rect 345782 516618 345866 516854
rect 346102 516618 379546 516854
rect 379782 516618 379866 516854
rect 380102 516618 413546 516854
rect 413782 516618 413866 516854
rect 414102 516618 447546 516854
rect 447782 516618 447866 516854
rect 448102 516618 481546 516854
rect 481782 516618 481866 516854
rect 482102 516618 515546 516854
rect 515782 516618 515866 516854
rect 516102 516618 549546 516854
rect 549782 516618 549866 516854
rect 550102 516618 586302 516854
rect 586538 516618 586622 516854
rect 586858 516618 592650 516854
rect -8726 516586 592650 516618
rect -8726 513454 592650 513486
rect -8726 513218 -1974 513454
rect -1738 513218 -1654 513454
rect -1418 513218 1826 513454
rect 2062 513218 2146 513454
rect 2382 513218 35826 513454
rect 36062 513218 36146 513454
rect 36382 513218 69826 513454
rect 70062 513218 70146 513454
rect 70382 513218 103826 513454
rect 104062 513218 104146 513454
rect 104382 513218 137826 513454
rect 138062 513218 138146 513454
rect 138382 513218 171826 513454
rect 172062 513218 172146 513454
rect 172382 513218 205826 513454
rect 206062 513218 206146 513454
rect 206382 513218 239826 513454
rect 240062 513218 240146 513454
rect 240382 513218 273826 513454
rect 274062 513218 274146 513454
rect 274382 513218 307826 513454
rect 308062 513218 308146 513454
rect 308382 513218 341826 513454
rect 342062 513218 342146 513454
rect 342382 513218 375826 513454
rect 376062 513218 376146 513454
rect 376382 513218 409826 513454
rect 410062 513218 410146 513454
rect 410382 513218 443826 513454
rect 444062 513218 444146 513454
rect 444382 513218 477826 513454
rect 478062 513218 478146 513454
rect 478382 513218 511826 513454
rect 512062 513218 512146 513454
rect 512382 513218 545826 513454
rect 546062 513218 546146 513454
rect 546382 513218 579826 513454
rect 580062 513218 580146 513454
rect 580382 513218 585342 513454
rect 585578 513218 585662 513454
rect 585898 513218 592650 513454
rect -8726 513134 592650 513218
rect -8726 512898 -1974 513134
rect -1738 512898 -1654 513134
rect -1418 512898 1826 513134
rect 2062 512898 2146 513134
rect 2382 512898 35826 513134
rect 36062 512898 36146 513134
rect 36382 512898 69826 513134
rect 70062 512898 70146 513134
rect 70382 512898 103826 513134
rect 104062 512898 104146 513134
rect 104382 512898 137826 513134
rect 138062 512898 138146 513134
rect 138382 512898 171826 513134
rect 172062 512898 172146 513134
rect 172382 512898 205826 513134
rect 206062 512898 206146 513134
rect 206382 512898 239826 513134
rect 240062 512898 240146 513134
rect 240382 512898 273826 513134
rect 274062 512898 274146 513134
rect 274382 512898 307826 513134
rect 308062 512898 308146 513134
rect 308382 512898 341826 513134
rect 342062 512898 342146 513134
rect 342382 512898 375826 513134
rect 376062 512898 376146 513134
rect 376382 512898 409826 513134
rect 410062 512898 410146 513134
rect 410382 512898 443826 513134
rect 444062 512898 444146 513134
rect 444382 512898 477826 513134
rect 478062 512898 478146 513134
rect 478382 512898 511826 513134
rect 512062 512898 512146 513134
rect 512382 512898 545826 513134
rect 546062 512898 546146 513134
rect 546382 512898 579826 513134
rect 580062 512898 580146 513134
rect 580382 512898 585342 513134
rect 585578 512898 585662 513134
rect 585898 512898 592650 513134
rect -8726 512866 592650 512898
rect -8726 505494 592650 505526
rect -8726 505258 -8694 505494
rect -8458 505258 -8374 505494
rect -8138 505258 27866 505494
rect 28102 505258 28186 505494
rect 28422 505258 61866 505494
rect 62102 505258 62186 505494
rect 62422 505258 95866 505494
rect 96102 505258 96186 505494
rect 96422 505258 129866 505494
rect 130102 505258 130186 505494
rect 130422 505258 163866 505494
rect 164102 505258 164186 505494
rect 164422 505258 197866 505494
rect 198102 505258 198186 505494
rect 198422 505258 231866 505494
rect 232102 505258 232186 505494
rect 232422 505258 265866 505494
rect 266102 505258 266186 505494
rect 266422 505258 299866 505494
rect 300102 505258 300186 505494
rect 300422 505258 333866 505494
rect 334102 505258 334186 505494
rect 334422 505258 367866 505494
rect 368102 505258 368186 505494
rect 368422 505258 401866 505494
rect 402102 505258 402186 505494
rect 402422 505258 435866 505494
rect 436102 505258 436186 505494
rect 436422 505258 469866 505494
rect 470102 505258 470186 505494
rect 470422 505258 503866 505494
rect 504102 505258 504186 505494
rect 504422 505258 537866 505494
rect 538102 505258 538186 505494
rect 538422 505258 571866 505494
rect 572102 505258 572186 505494
rect 572422 505258 592062 505494
rect 592298 505258 592382 505494
rect 592618 505258 592650 505494
rect -8726 505174 592650 505258
rect -8726 504938 -8694 505174
rect -8458 504938 -8374 505174
rect -8138 504938 27866 505174
rect 28102 504938 28186 505174
rect 28422 504938 61866 505174
rect 62102 504938 62186 505174
rect 62422 504938 95866 505174
rect 96102 504938 96186 505174
rect 96422 504938 129866 505174
rect 130102 504938 130186 505174
rect 130422 504938 163866 505174
rect 164102 504938 164186 505174
rect 164422 504938 197866 505174
rect 198102 504938 198186 505174
rect 198422 504938 231866 505174
rect 232102 504938 232186 505174
rect 232422 504938 265866 505174
rect 266102 504938 266186 505174
rect 266422 504938 299866 505174
rect 300102 504938 300186 505174
rect 300422 504938 333866 505174
rect 334102 504938 334186 505174
rect 334422 504938 367866 505174
rect 368102 504938 368186 505174
rect 368422 504938 401866 505174
rect 402102 504938 402186 505174
rect 402422 504938 435866 505174
rect 436102 504938 436186 505174
rect 436422 504938 469866 505174
rect 470102 504938 470186 505174
rect 470422 504938 503866 505174
rect 504102 504938 504186 505174
rect 504422 504938 537866 505174
rect 538102 504938 538186 505174
rect 538422 504938 571866 505174
rect 572102 504938 572186 505174
rect 572422 504938 592062 505174
rect 592298 504938 592382 505174
rect 592618 504938 592650 505174
rect -8726 504906 592650 504938
rect -8726 501774 592650 501806
rect -8726 501538 -7734 501774
rect -7498 501538 -7414 501774
rect -7178 501538 24146 501774
rect 24382 501538 24466 501774
rect 24702 501538 58146 501774
rect 58382 501538 58466 501774
rect 58702 501538 92146 501774
rect 92382 501538 92466 501774
rect 92702 501538 126146 501774
rect 126382 501538 126466 501774
rect 126702 501538 160146 501774
rect 160382 501538 160466 501774
rect 160702 501538 194146 501774
rect 194382 501538 194466 501774
rect 194702 501538 228146 501774
rect 228382 501538 228466 501774
rect 228702 501538 262146 501774
rect 262382 501538 262466 501774
rect 262702 501538 296146 501774
rect 296382 501538 296466 501774
rect 296702 501538 330146 501774
rect 330382 501538 330466 501774
rect 330702 501538 364146 501774
rect 364382 501538 364466 501774
rect 364702 501538 398146 501774
rect 398382 501538 398466 501774
rect 398702 501538 432146 501774
rect 432382 501538 432466 501774
rect 432702 501538 466146 501774
rect 466382 501538 466466 501774
rect 466702 501538 500146 501774
rect 500382 501538 500466 501774
rect 500702 501538 534146 501774
rect 534382 501538 534466 501774
rect 534702 501538 568146 501774
rect 568382 501538 568466 501774
rect 568702 501538 591102 501774
rect 591338 501538 591422 501774
rect 591658 501538 592650 501774
rect -8726 501454 592650 501538
rect -8726 501218 -7734 501454
rect -7498 501218 -7414 501454
rect -7178 501218 24146 501454
rect 24382 501218 24466 501454
rect 24702 501218 58146 501454
rect 58382 501218 58466 501454
rect 58702 501218 92146 501454
rect 92382 501218 92466 501454
rect 92702 501218 126146 501454
rect 126382 501218 126466 501454
rect 126702 501218 160146 501454
rect 160382 501218 160466 501454
rect 160702 501218 194146 501454
rect 194382 501218 194466 501454
rect 194702 501218 228146 501454
rect 228382 501218 228466 501454
rect 228702 501218 262146 501454
rect 262382 501218 262466 501454
rect 262702 501218 296146 501454
rect 296382 501218 296466 501454
rect 296702 501218 330146 501454
rect 330382 501218 330466 501454
rect 330702 501218 364146 501454
rect 364382 501218 364466 501454
rect 364702 501218 398146 501454
rect 398382 501218 398466 501454
rect 398702 501218 432146 501454
rect 432382 501218 432466 501454
rect 432702 501218 466146 501454
rect 466382 501218 466466 501454
rect 466702 501218 500146 501454
rect 500382 501218 500466 501454
rect 500702 501218 534146 501454
rect 534382 501218 534466 501454
rect 534702 501218 568146 501454
rect 568382 501218 568466 501454
rect 568702 501218 591102 501454
rect 591338 501218 591422 501454
rect 591658 501218 592650 501454
rect -8726 501186 592650 501218
rect -8726 498054 592650 498086
rect -8726 497818 -6774 498054
rect -6538 497818 -6454 498054
rect -6218 497818 20426 498054
rect 20662 497818 20746 498054
rect 20982 497818 54426 498054
rect 54662 497818 54746 498054
rect 54982 497818 88426 498054
rect 88662 497818 88746 498054
rect 88982 497818 122426 498054
rect 122662 497818 122746 498054
rect 122982 497818 156426 498054
rect 156662 497818 156746 498054
rect 156982 497818 190426 498054
rect 190662 497818 190746 498054
rect 190982 497818 224426 498054
rect 224662 497818 224746 498054
rect 224982 497818 258426 498054
rect 258662 497818 258746 498054
rect 258982 497818 292426 498054
rect 292662 497818 292746 498054
rect 292982 497818 326426 498054
rect 326662 497818 326746 498054
rect 326982 497818 360426 498054
rect 360662 497818 360746 498054
rect 360982 497818 394426 498054
rect 394662 497818 394746 498054
rect 394982 497818 428426 498054
rect 428662 497818 428746 498054
rect 428982 497818 462426 498054
rect 462662 497818 462746 498054
rect 462982 497818 496426 498054
rect 496662 497818 496746 498054
rect 496982 497818 530426 498054
rect 530662 497818 530746 498054
rect 530982 497818 564426 498054
rect 564662 497818 564746 498054
rect 564982 497818 590142 498054
rect 590378 497818 590462 498054
rect 590698 497818 592650 498054
rect -8726 497734 592650 497818
rect -8726 497498 -6774 497734
rect -6538 497498 -6454 497734
rect -6218 497498 20426 497734
rect 20662 497498 20746 497734
rect 20982 497498 54426 497734
rect 54662 497498 54746 497734
rect 54982 497498 88426 497734
rect 88662 497498 88746 497734
rect 88982 497498 122426 497734
rect 122662 497498 122746 497734
rect 122982 497498 156426 497734
rect 156662 497498 156746 497734
rect 156982 497498 190426 497734
rect 190662 497498 190746 497734
rect 190982 497498 224426 497734
rect 224662 497498 224746 497734
rect 224982 497498 258426 497734
rect 258662 497498 258746 497734
rect 258982 497498 292426 497734
rect 292662 497498 292746 497734
rect 292982 497498 326426 497734
rect 326662 497498 326746 497734
rect 326982 497498 360426 497734
rect 360662 497498 360746 497734
rect 360982 497498 394426 497734
rect 394662 497498 394746 497734
rect 394982 497498 428426 497734
rect 428662 497498 428746 497734
rect 428982 497498 462426 497734
rect 462662 497498 462746 497734
rect 462982 497498 496426 497734
rect 496662 497498 496746 497734
rect 496982 497498 530426 497734
rect 530662 497498 530746 497734
rect 530982 497498 564426 497734
rect 564662 497498 564746 497734
rect 564982 497498 590142 497734
rect 590378 497498 590462 497734
rect 590698 497498 592650 497734
rect -8726 497466 592650 497498
rect -8726 494334 592650 494366
rect -8726 494098 -5814 494334
rect -5578 494098 -5494 494334
rect -5258 494098 16706 494334
rect 16942 494098 17026 494334
rect 17262 494098 50706 494334
rect 50942 494098 51026 494334
rect 51262 494098 84706 494334
rect 84942 494098 85026 494334
rect 85262 494098 118706 494334
rect 118942 494098 119026 494334
rect 119262 494098 152706 494334
rect 152942 494098 153026 494334
rect 153262 494098 186706 494334
rect 186942 494098 187026 494334
rect 187262 494098 220706 494334
rect 220942 494098 221026 494334
rect 221262 494098 254706 494334
rect 254942 494098 255026 494334
rect 255262 494098 288706 494334
rect 288942 494098 289026 494334
rect 289262 494098 322706 494334
rect 322942 494098 323026 494334
rect 323262 494098 356706 494334
rect 356942 494098 357026 494334
rect 357262 494098 390706 494334
rect 390942 494098 391026 494334
rect 391262 494098 424706 494334
rect 424942 494098 425026 494334
rect 425262 494098 458706 494334
rect 458942 494098 459026 494334
rect 459262 494098 492706 494334
rect 492942 494098 493026 494334
rect 493262 494098 526706 494334
rect 526942 494098 527026 494334
rect 527262 494098 560706 494334
rect 560942 494098 561026 494334
rect 561262 494098 589182 494334
rect 589418 494098 589502 494334
rect 589738 494098 592650 494334
rect -8726 494014 592650 494098
rect -8726 493778 -5814 494014
rect -5578 493778 -5494 494014
rect -5258 493778 16706 494014
rect 16942 493778 17026 494014
rect 17262 493778 50706 494014
rect 50942 493778 51026 494014
rect 51262 493778 84706 494014
rect 84942 493778 85026 494014
rect 85262 493778 118706 494014
rect 118942 493778 119026 494014
rect 119262 493778 152706 494014
rect 152942 493778 153026 494014
rect 153262 493778 186706 494014
rect 186942 493778 187026 494014
rect 187262 493778 220706 494014
rect 220942 493778 221026 494014
rect 221262 493778 254706 494014
rect 254942 493778 255026 494014
rect 255262 493778 288706 494014
rect 288942 493778 289026 494014
rect 289262 493778 322706 494014
rect 322942 493778 323026 494014
rect 323262 493778 356706 494014
rect 356942 493778 357026 494014
rect 357262 493778 390706 494014
rect 390942 493778 391026 494014
rect 391262 493778 424706 494014
rect 424942 493778 425026 494014
rect 425262 493778 458706 494014
rect 458942 493778 459026 494014
rect 459262 493778 492706 494014
rect 492942 493778 493026 494014
rect 493262 493778 526706 494014
rect 526942 493778 527026 494014
rect 527262 493778 560706 494014
rect 560942 493778 561026 494014
rect 561262 493778 589182 494014
rect 589418 493778 589502 494014
rect 589738 493778 592650 494014
rect -8726 493746 592650 493778
rect -8726 490614 592650 490646
rect -8726 490378 -4854 490614
rect -4618 490378 -4534 490614
rect -4298 490378 12986 490614
rect 13222 490378 13306 490614
rect 13542 490378 46986 490614
rect 47222 490378 47306 490614
rect 47542 490378 80986 490614
rect 81222 490378 81306 490614
rect 81542 490378 114986 490614
rect 115222 490378 115306 490614
rect 115542 490378 148986 490614
rect 149222 490378 149306 490614
rect 149542 490378 182986 490614
rect 183222 490378 183306 490614
rect 183542 490378 216986 490614
rect 217222 490378 217306 490614
rect 217542 490378 250986 490614
rect 251222 490378 251306 490614
rect 251542 490378 284986 490614
rect 285222 490378 285306 490614
rect 285542 490378 318986 490614
rect 319222 490378 319306 490614
rect 319542 490378 352986 490614
rect 353222 490378 353306 490614
rect 353542 490378 386986 490614
rect 387222 490378 387306 490614
rect 387542 490378 420986 490614
rect 421222 490378 421306 490614
rect 421542 490378 454986 490614
rect 455222 490378 455306 490614
rect 455542 490378 488986 490614
rect 489222 490378 489306 490614
rect 489542 490378 522986 490614
rect 523222 490378 523306 490614
rect 523542 490378 556986 490614
rect 557222 490378 557306 490614
rect 557542 490378 588222 490614
rect 588458 490378 588542 490614
rect 588778 490378 592650 490614
rect -8726 490294 592650 490378
rect -8726 490058 -4854 490294
rect -4618 490058 -4534 490294
rect -4298 490058 12986 490294
rect 13222 490058 13306 490294
rect 13542 490058 46986 490294
rect 47222 490058 47306 490294
rect 47542 490058 80986 490294
rect 81222 490058 81306 490294
rect 81542 490058 114986 490294
rect 115222 490058 115306 490294
rect 115542 490058 148986 490294
rect 149222 490058 149306 490294
rect 149542 490058 182986 490294
rect 183222 490058 183306 490294
rect 183542 490058 216986 490294
rect 217222 490058 217306 490294
rect 217542 490058 250986 490294
rect 251222 490058 251306 490294
rect 251542 490058 284986 490294
rect 285222 490058 285306 490294
rect 285542 490058 318986 490294
rect 319222 490058 319306 490294
rect 319542 490058 352986 490294
rect 353222 490058 353306 490294
rect 353542 490058 386986 490294
rect 387222 490058 387306 490294
rect 387542 490058 420986 490294
rect 421222 490058 421306 490294
rect 421542 490058 454986 490294
rect 455222 490058 455306 490294
rect 455542 490058 488986 490294
rect 489222 490058 489306 490294
rect 489542 490058 522986 490294
rect 523222 490058 523306 490294
rect 523542 490058 556986 490294
rect 557222 490058 557306 490294
rect 557542 490058 588222 490294
rect 588458 490058 588542 490294
rect 588778 490058 592650 490294
rect -8726 490026 592650 490058
rect -8726 486894 592650 486926
rect -8726 486658 -3894 486894
rect -3658 486658 -3574 486894
rect -3338 486658 9266 486894
rect 9502 486658 9586 486894
rect 9822 486658 43266 486894
rect 43502 486658 43586 486894
rect 43822 486658 77266 486894
rect 77502 486658 77586 486894
rect 77822 486658 111266 486894
rect 111502 486658 111586 486894
rect 111822 486658 145266 486894
rect 145502 486658 145586 486894
rect 145822 486658 179266 486894
rect 179502 486658 179586 486894
rect 179822 486658 213266 486894
rect 213502 486658 213586 486894
rect 213822 486658 247266 486894
rect 247502 486658 247586 486894
rect 247822 486658 281266 486894
rect 281502 486658 281586 486894
rect 281822 486658 315266 486894
rect 315502 486658 315586 486894
rect 315822 486658 349266 486894
rect 349502 486658 349586 486894
rect 349822 486658 383266 486894
rect 383502 486658 383586 486894
rect 383822 486658 417266 486894
rect 417502 486658 417586 486894
rect 417822 486658 451266 486894
rect 451502 486658 451586 486894
rect 451822 486658 485266 486894
rect 485502 486658 485586 486894
rect 485822 486658 519266 486894
rect 519502 486658 519586 486894
rect 519822 486658 553266 486894
rect 553502 486658 553586 486894
rect 553822 486658 587262 486894
rect 587498 486658 587582 486894
rect 587818 486658 592650 486894
rect -8726 486574 592650 486658
rect -8726 486338 -3894 486574
rect -3658 486338 -3574 486574
rect -3338 486338 9266 486574
rect 9502 486338 9586 486574
rect 9822 486338 43266 486574
rect 43502 486338 43586 486574
rect 43822 486338 77266 486574
rect 77502 486338 77586 486574
rect 77822 486338 111266 486574
rect 111502 486338 111586 486574
rect 111822 486338 145266 486574
rect 145502 486338 145586 486574
rect 145822 486338 179266 486574
rect 179502 486338 179586 486574
rect 179822 486338 213266 486574
rect 213502 486338 213586 486574
rect 213822 486338 247266 486574
rect 247502 486338 247586 486574
rect 247822 486338 281266 486574
rect 281502 486338 281586 486574
rect 281822 486338 315266 486574
rect 315502 486338 315586 486574
rect 315822 486338 349266 486574
rect 349502 486338 349586 486574
rect 349822 486338 383266 486574
rect 383502 486338 383586 486574
rect 383822 486338 417266 486574
rect 417502 486338 417586 486574
rect 417822 486338 451266 486574
rect 451502 486338 451586 486574
rect 451822 486338 485266 486574
rect 485502 486338 485586 486574
rect 485822 486338 519266 486574
rect 519502 486338 519586 486574
rect 519822 486338 553266 486574
rect 553502 486338 553586 486574
rect 553822 486338 587262 486574
rect 587498 486338 587582 486574
rect 587818 486338 592650 486574
rect -8726 486306 592650 486338
rect -8726 483174 592650 483206
rect -8726 482938 -2934 483174
rect -2698 482938 -2614 483174
rect -2378 482938 5546 483174
rect 5782 482938 5866 483174
rect 6102 482938 39546 483174
rect 39782 482938 39866 483174
rect 40102 482938 73546 483174
rect 73782 482938 73866 483174
rect 74102 482938 107546 483174
rect 107782 482938 107866 483174
rect 108102 482938 141546 483174
rect 141782 482938 141866 483174
rect 142102 482938 175546 483174
rect 175782 482938 175866 483174
rect 176102 482938 209546 483174
rect 209782 482938 209866 483174
rect 210102 482938 243546 483174
rect 243782 482938 243866 483174
rect 244102 482938 277546 483174
rect 277782 482938 277866 483174
rect 278102 482938 311546 483174
rect 311782 482938 311866 483174
rect 312102 482938 345546 483174
rect 345782 482938 345866 483174
rect 346102 482938 379546 483174
rect 379782 482938 379866 483174
rect 380102 482938 413546 483174
rect 413782 482938 413866 483174
rect 414102 482938 447546 483174
rect 447782 482938 447866 483174
rect 448102 482938 481546 483174
rect 481782 482938 481866 483174
rect 482102 482938 515546 483174
rect 515782 482938 515866 483174
rect 516102 482938 549546 483174
rect 549782 482938 549866 483174
rect 550102 482938 586302 483174
rect 586538 482938 586622 483174
rect 586858 482938 592650 483174
rect -8726 482854 592650 482938
rect -8726 482618 -2934 482854
rect -2698 482618 -2614 482854
rect -2378 482618 5546 482854
rect 5782 482618 5866 482854
rect 6102 482618 39546 482854
rect 39782 482618 39866 482854
rect 40102 482618 73546 482854
rect 73782 482618 73866 482854
rect 74102 482618 107546 482854
rect 107782 482618 107866 482854
rect 108102 482618 141546 482854
rect 141782 482618 141866 482854
rect 142102 482618 175546 482854
rect 175782 482618 175866 482854
rect 176102 482618 209546 482854
rect 209782 482618 209866 482854
rect 210102 482618 243546 482854
rect 243782 482618 243866 482854
rect 244102 482618 277546 482854
rect 277782 482618 277866 482854
rect 278102 482618 311546 482854
rect 311782 482618 311866 482854
rect 312102 482618 345546 482854
rect 345782 482618 345866 482854
rect 346102 482618 379546 482854
rect 379782 482618 379866 482854
rect 380102 482618 413546 482854
rect 413782 482618 413866 482854
rect 414102 482618 447546 482854
rect 447782 482618 447866 482854
rect 448102 482618 481546 482854
rect 481782 482618 481866 482854
rect 482102 482618 515546 482854
rect 515782 482618 515866 482854
rect 516102 482618 549546 482854
rect 549782 482618 549866 482854
rect 550102 482618 586302 482854
rect 586538 482618 586622 482854
rect 586858 482618 592650 482854
rect -8726 482586 592650 482618
rect -8726 479454 592650 479486
rect -8726 479218 -1974 479454
rect -1738 479218 -1654 479454
rect -1418 479218 1826 479454
rect 2062 479218 2146 479454
rect 2382 479218 35826 479454
rect 36062 479218 36146 479454
rect 36382 479218 69826 479454
rect 70062 479218 70146 479454
rect 70382 479218 103826 479454
rect 104062 479218 104146 479454
rect 104382 479218 137826 479454
rect 138062 479218 138146 479454
rect 138382 479218 171826 479454
rect 172062 479218 172146 479454
rect 172382 479218 205826 479454
rect 206062 479218 206146 479454
rect 206382 479218 239826 479454
rect 240062 479218 240146 479454
rect 240382 479218 273826 479454
rect 274062 479218 274146 479454
rect 274382 479218 307826 479454
rect 308062 479218 308146 479454
rect 308382 479218 341826 479454
rect 342062 479218 342146 479454
rect 342382 479218 375826 479454
rect 376062 479218 376146 479454
rect 376382 479218 409826 479454
rect 410062 479218 410146 479454
rect 410382 479218 443826 479454
rect 444062 479218 444146 479454
rect 444382 479218 477826 479454
rect 478062 479218 478146 479454
rect 478382 479218 511826 479454
rect 512062 479218 512146 479454
rect 512382 479218 545826 479454
rect 546062 479218 546146 479454
rect 546382 479218 579826 479454
rect 580062 479218 580146 479454
rect 580382 479218 585342 479454
rect 585578 479218 585662 479454
rect 585898 479218 592650 479454
rect -8726 479134 592650 479218
rect -8726 478898 -1974 479134
rect -1738 478898 -1654 479134
rect -1418 478898 1826 479134
rect 2062 478898 2146 479134
rect 2382 478898 35826 479134
rect 36062 478898 36146 479134
rect 36382 478898 69826 479134
rect 70062 478898 70146 479134
rect 70382 478898 103826 479134
rect 104062 478898 104146 479134
rect 104382 478898 137826 479134
rect 138062 478898 138146 479134
rect 138382 478898 171826 479134
rect 172062 478898 172146 479134
rect 172382 478898 205826 479134
rect 206062 478898 206146 479134
rect 206382 478898 239826 479134
rect 240062 478898 240146 479134
rect 240382 478898 273826 479134
rect 274062 478898 274146 479134
rect 274382 478898 307826 479134
rect 308062 478898 308146 479134
rect 308382 478898 341826 479134
rect 342062 478898 342146 479134
rect 342382 478898 375826 479134
rect 376062 478898 376146 479134
rect 376382 478898 409826 479134
rect 410062 478898 410146 479134
rect 410382 478898 443826 479134
rect 444062 478898 444146 479134
rect 444382 478898 477826 479134
rect 478062 478898 478146 479134
rect 478382 478898 511826 479134
rect 512062 478898 512146 479134
rect 512382 478898 545826 479134
rect 546062 478898 546146 479134
rect 546382 478898 579826 479134
rect 580062 478898 580146 479134
rect 580382 478898 585342 479134
rect 585578 478898 585662 479134
rect 585898 478898 592650 479134
rect -8726 478866 592650 478898
rect -8726 471494 592650 471526
rect -8726 471258 -8694 471494
rect -8458 471258 -8374 471494
rect -8138 471258 27866 471494
rect 28102 471258 28186 471494
rect 28422 471258 61866 471494
rect 62102 471258 62186 471494
rect 62422 471258 95866 471494
rect 96102 471258 96186 471494
rect 96422 471258 129866 471494
rect 130102 471258 130186 471494
rect 130422 471258 163866 471494
rect 164102 471258 164186 471494
rect 164422 471258 197866 471494
rect 198102 471258 198186 471494
rect 198422 471258 231866 471494
rect 232102 471258 232186 471494
rect 232422 471258 265866 471494
rect 266102 471258 266186 471494
rect 266422 471258 299866 471494
rect 300102 471258 300186 471494
rect 300422 471258 333866 471494
rect 334102 471258 334186 471494
rect 334422 471258 367866 471494
rect 368102 471258 368186 471494
rect 368422 471258 401866 471494
rect 402102 471258 402186 471494
rect 402422 471258 435866 471494
rect 436102 471258 436186 471494
rect 436422 471258 469866 471494
rect 470102 471258 470186 471494
rect 470422 471258 503866 471494
rect 504102 471258 504186 471494
rect 504422 471258 537866 471494
rect 538102 471258 538186 471494
rect 538422 471258 571866 471494
rect 572102 471258 572186 471494
rect 572422 471258 592062 471494
rect 592298 471258 592382 471494
rect 592618 471258 592650 471494
rect -8726 471174 592650 471258
rect -8726 470938 -8694 471174
rect -8458 470938 -8374 471174
rect -8138 470938 27866 471174
rect 28102 470938 28186 471174
rect 28422 470938 61866 471174
rect 62102 470938 62186 471174
rect 62422 470938 95866 471174
rect 96102 470938 96186 471174
rect 96422 470938 129866 471174
rect 130102 470938 130186 471174
rect 130422 470938 163866 471174
rect 164102 470938 164186 471174
rect 164422 470938 197866 471174
rect 198102 470938 198186 471174
rect 198422 470938 231866 471174
rect 232102 470938 232186 471174
rect 232422 470938 265866 471174
rect 266102 470938 266186 471174
rect 266422 470938 299866 471174
rect 300102 470938 300186 471174
rect 300422 470938 333866 471174
rect 334102 470938 334186 471174
rect 334422 470938 367866 471174
rect 368102 470938 368186 471174
rect 368422 470938 401866 471174
rect 402102 470938 402186 471174
rect 402422 470938 435866 471174
rect 436102 470938 436186 471174
rect 436422 470938 469866 471174
rect 470102 470938 470186 471174
rect 470422 470938 503866 471174
rect 504102 470938 504186 471174
rect 504422 470938 537866 471174
rect 538102 470938 538186 471174
rect 538422 470938 571866 471174
rect 572102 470938 572186 471174
rect 572422 470938 592062 471174
rect 592298 470938 592382 471174
rect 592618 470938 592650 471174
rect -8726 470906 592650 470938
rect -8726 467774 592650 467806
rect -8726 467538 -7734 467774
rect -7498 467538 -7414 467774
rect -7178 467538 24146 467774
rect 24382 467538 24466 467774
rect 24702 467538 58146 467774
rect 58382 467538 58466 467774
rect 58702 467538 92146 467774
rect 92382 467538 92466 467774
rect 92702 467538 126146 467774
rect 126382 467538 126466 467774
rect 126702 467538 160146 467774
rect 160382 467538 160466 467774
rect 160702 467538 194146 467774
rect 194382 467538 194466 467774
rect 194702 467538 228146 467774
rect 228382 467538 228466 467774
rect 228702 467538 262146 467774
rect 262382 467538 262466 467774
rect 262702 467538 296146 467774
rect 296382 467538 296466 467774
rect 296702 467538 330146 467774
rect 330382 467538 330466 467774
rect 330702 467538 364146 467774
rect 364382 467538 364466 467774
rect 364702 467538 398146 467774
rect 398382 467538 398466 467774
rect 398702 467538 432146 467774
rect 432382 467538 432466 467774
rect 432702 467538 466146 467774
rect 466382 467538 466466 467774
rect 466702 467538 500146 467774
rect 500382 467538 500466 467774
rect 500702 467538 534146 467774
rect 534382 467538 534466 467774
rect 534702 467538 568146 467774
rect 568382 467538 568466 467774
rect 568702 467538 591102 467774
rect 591338 467538 591422 467774
rect 591658 467538 592650 467774
rect -8726 467454 592650 467538
rect -8726 467218 -7734 467454
rect -7498 467218 -7414 467454
rect -7178 467218 24146 467454
rect 24382 467218 24466 467454
rect 24702 467218 58146 467454
rect 58382 467218 58466 467454
rect 58702 467218 92146 467454
rect 92382 467218 92466 467454
rect 92702 467218 126146 467454
rect 126382 467218 126466 467454
rect 126702 467218 160146 467454
rect 160382 467218 160466 467454
rect 160702 467218 194146 467454
rect 194382 467218 194466 467454
rect 194702 467218 228146 467454
rect 228382 467218 228466 467454
rect 228702 467218 262146 467454
rect 262382 467218 262466 467454
rect 262702 467218 296146 467454
rect 296382 467218 296466 467454
rect 296702 467218 330146 467454
rect 330382 467218 330466 467454
rect 330702 467218 364146 467454
rect 364382 467218 364466 467454
rect 364702 467218 398146 467454
rect 398382 467218 398466 467454
rect 398702 467218 432146 467454
rect 432382 467218 432466 467454
rect 432702 467218 466146 467454
rect 466382 467218 466466 467454
rect 466702 467218 500146 467454
rect 500382 467218 500466 467454
rect 500702 467218 534146 467454
rect 534382 467218 534466 467454
rect 534702 467218 568146 467454
rect 568382 467218 568466 467454
rect 568702 467218 591102 467454
rect 591338 467218 591422 467454
rect 591658 467218 592650 467454
rect -8726 467186 592650 467218
rect -8726 464054 592650 464086
rect -8726 463818 -6774 464054
rect -6538 463818 -6454 464054
rect -6218 463818 20426 464054
rect 20662 463818 20746 464054
rect 20982 463818 54426 464054
rect 54662 463818 54746 464054
rect 54982 463818 88426 464054
rect 88662 463818 88746 464054
rect 88982 463818 122426 464054
rect 122662 463818 122746 464054
rect 122982 463818 156426 464054
rect 156662 463818 156746 464054
rect 156982 463818 190426 464054
rect 190662 463818 190746 464054
rect 190982 463818 224426 464054
rect 224662 463818 224746 464054
rect 224982 463818 258426 464054
rect 258662 463818 258746 464054
rect 258982 463818 292426 464054
rect 292662 463818 292746 464054
rect 292982 463818 326426 464054
rect 326662 463818 326746 464054
rect 326982 463818 360426 464054
rect 360662 463818 360746 464054
rect 360982 463818 394426 464054
rect 394662 463818 394746 464054
rect 394982 463818 428426 464054
rect 428662 463818 428746 464054
rect 428982 463818 462426 464054
rect 462662 463818 462746 464054
rect 462982 463818 496426 464054
rect 496662 463818 496746 464054
rect 496982 463818 530426 464054
rect 530662 463818 530746 464054
rect 530982 463818 564426 464054
rect 564662 463818 564746 464054
rect 564982 463818 590142 464054
rect 590378 463818 590462 464054
rect 590698 463818 592650 464054
rect -8726 463734 592650 463818
rect -8726 463498 -6774 463734
rect -6538 463498 -6454 463734
rect -6218 463498 20426 463734
rect 20662 463498 20746 463734
rect 20982 463498 54426 463734
rect 54662 463498 54746 463734
rect 54982 463498 88426 463734
rect 88662 463498 88746 463734
rect 88982 463498 122426 463734
rect 122662 463498 122746 463734
rect 122982 463498 156426 463734
rect 156662 463498 156746 463734
rect 156982 463498 190426 463734
rect 190662 463498 190746 463734
rect 190982 463498 224426 463734
rect 224662 463498 224746 463734
rect 224982 463498 258426 463734
rect 258662 463498 258746 463734
rect 258982 463498 292426 463734
rect 292662 463498 292746 463734
rect 292982 463498 326426 463734
rect 326662 463498 326746 463734
rect 326982 463498 360426 463734
rect 360662 463498 360746 463734
rect 360982 463498 394426 463734
rect 394662 463498 394746 463734
rect 394982 463498 428426 463734
rect 428662 463498 428746 463734
rect 428982 463498 462426 463734
rect 462662 463498 462746 463734
rect 462982 463498 496426 463734
rect 496662 463498 496746 463734
rect 496982 463498 530426 463734
rect 530662 463498 530746 463734
rect 530982 463498 564426 463734
rect 564662 463498 564746 463734
rect 564982 463498 590142 463734
rect 590378 463498 590462 463734
rect 590698 463498 592650 463734
rect -8726 463466 592650 463498
rect -8726 460334 592650 460366
rect -8726 460098 -5814 460334
rect -5578 460098 -5494 460334
rect -5258 460098 16706 460334
rect 16942 460098 17026 460334
rect 17262 460098 50706 460334
rect 50942 460098 51026 460334
rect 51262 460098 84706 460334
rect 84942 460098 85026 460334
rect 85262 460098 118706 460334
rect 118942 460098 119026 460334
rect 119262 460098 152706 460334
rect 152942 460098 153026 460334
rect 153262 460098 186706 460334
rect 186942 460098 187026 460334
rect 187262 460098 220706 460334
rect 220942 460098 221026 460334
rect 221262 460098 254706 460334
rect 254942 460098 255026 460334
rect 255262 460098 288706 460334
rect 288942 460098 289026 460334
rect 289262 460098 322706 460334
rect 322942 460098 323026 460334
rect 323262 460098 356706 460334
rect 356942 460098 357026 460334
rect 357262 460098 390706 460334
rect 390942 460098 391026 460334
rect 391262 460098 424706 460334
rect 424942 460098 425026 460334
rect 425262 460098 458706 460334
rect 458942 460098 459026 460334
rect 459262 460098 492706 460334
rect 492942 460098 493026 460334
rect 493262 460098 526706 460334
rect 526942 460098 527026 460334
rect 527262 460098 560706 460334
rect 560942 460098 561026 460334
rect 561262 460098 589182 460334
rect 589418 460098 589502 460334
rect 589738 460098 592650 460334
rect -8726 460014 592650 460098
rect -8726 459778 -5814 460014
rect -5578 459778 -5494 460014
rect -5258 459778 16706 460014
rect 16942 459778 17026 460014
rect 17262 459778 50706 460014
rect 50942 459778 51026 460014
rect 51262 459778 84706 460014
rect 84942 459778 85026 460014
rect 85262 459778 118706 460014
rect 118942 459778 119026 460014
rect 119262 459778 152706 460014
rect 152942 459778 153026 460014
rect 153262 459778 186706 460014
rect 186942 459778 187026 460014
rect 187262 459778 220706 460014
rect 220942 459778 221026 460014
rect 221262 459778 254706 460014
rect 254942 459778 255026 460014
rect 255262 459778 288706 460014
rect 288942 459778 289026 460014
rect 289262 459778 322706 460014
rect 322942 459778 323026 460014
rect 323262 459778 356706 460014
rect 356942 459778 357026 460014
rect 357262 459778 390706 460014
rect 390942 459778 391026 460014
rect 391262 459778 424706 460014
rect 424942 459778 425026 460014
rect 425262 459778 458706 460014
rect 458942 459778 459026 460014
rect 459262 459778 492706 460014
rect 492942 459778 493026 460014
rect 493262 459778 526706 460014
rect 526942 459778 527026 460014
rect 527262 459778 560706 460014
rect 560942 459778 561026 460014
rect 561262 459778 589182 460014
rect 589418 459778 589502 460014
rect 589738 459778 592650 460014
rect -8726 459746 592650 459778
rect -8726 456614 592650 456646
rect -8726 456378 -4854 456614
rect -4618 456378 -4534 456614
rect -4298 456378 12986 456614
rect 13222 456378 13306 456614
rect 13542 456378 46986 456614
rect 47222 456378 47306 456614
rect 47542 456378 80986 456614
rect 81222 456378 81306 456614
rect 81542 456378 114986 456614
rect 115222 456378 115306 456614
rect 115542 456378 148986 456614
rect 149222 456378 149306 456614
rect 149542 456378 182986 456614
rect 183222 456378 183306 456614
rect 183542 456378 216986 456614
rect 217222 456378 217306 456614
rect 217542 456378 250986 456614
rect 251222 456378 251306 456614
rect 251542 456378 284986 456614
rect 285222 456378 285306 456614
rect 285542 456378 318986 456614
rect 319222 456378 319306 456614
rect 319542 456378 352986 456614
rect 353222 456378 353306 456614
rect 353542 456378 386986 456614
rect 387222 456378 387306 456614
rect 387542 456378 420986 456614
rect 421222 456378 421306 456614
rect 421542 456378 454986 456614
rect 455222 456378 455306 456614
rect 455542 456378 488986 456614
rect 489222 456378 489306 456614
rect 489542 456378 522986 456614
rect 523222 456378 523306 456614
rect 523542 456378 556986 456614
rect 557222 456378 557306 456614
rect 557542 456378 588222 456614
rect 588458 456378 588542 456614
rect 588778 456378 592650 456614
rect -8726 456294 592650 456378
rect -8726 456058 -4854 456294
rect -4618 456058 -4534 456294
rect -4298 456058 12986 456294
rect 13222 456058 13306 456294
rect 13542 456058 46986 456294
rect 47222 456058 47306 456294
rect 47542 456058 80986 456294
rect 81222 456058 81306 456294
rect 81542 456058 114986 456294
rect 115222 456058 115306 456294
rect 115542 456058 148986 456294
rect 149222 456058 149306 456294
rect 149542 456058 182986 456294
rect 183222 456058 183306 456294
rect 183542 456058 216986 456294
rect 217222 456058 217306 456294
rect 217542 456058 250986 456294
rect 251222 456058 251306 456294
rect 251542 456058 284986 456294
rect 285222 456058 285306 456294
rect 285542 456058 318986 456294
rect 319222 456058 319306 456294
rect 319542 456058 352986 456294
rect 353222 456058 353306 456294
rect 353542 456058 386986 456294
rect 387222 456058 387306 456294
rect 387542 456058 420986 456294
rect 421222 456058 421306 456294
rect 421542 456058 454986 456294
rect 455222 456058 455306 456294
rect 455542 456058 488986 456294
rect 489222 456058 489306 456294
rect 489542 456058 522986 456294
rect 523222 456058 523306 456294
rect 523542 456058 556986 456294
rect 557222 456058 557306 456294
rect 557542 456058 588222 456294
rect 588458 456058 588542 456294
rect 588778 456058 592650 456294
rect -8726 456026 592650 456058
rect -8726 452894 592650 452926
rect -8726 452658 -3894 452894
rect -3658 452658 -3574 452894
rect -3338 452658 9266 452894
rect 9502 452658 9586 452894
rect 9822 452658 43266 452894
rect 43502 452658 43586 452894
rect 43822 452658 77266 452894
rect 77502 452658 77586 452894
rect 77822 452658 111266 452894
rect 111502 452658 111586 452894
rect 111822 452658 145266 452894
rect 145502 452658 145586 452894
rect 145822 452658 179266 452894
rect 179502 452658 179586 452894
rect 179822 452658 213266 452894
rect 213502 452658 213586 452894
rect 213822 452658 247266 452894
rect 247502 452658 247586 452894
rect 247822 452658 281266 452894
rect 281502 452658 281586 452894
rect 281822 452658 315266 452894
rect 315502 452658 315586 452894
rect 315822 452658 349266 452894
rect 349502 452658 349586 452894
rect 349822 452658 383266 452894
rect 383502 452658 383586 452894
rect 383822 452658 417266 452894
rect 417502 452658 417586 452894
rect 417822 452658 451266 452894
rect 451502 452658 451586 452894
rect 451822 452658 485266 452894
rect 485502 452658 485586 452894
rect 485822 452658 519266 452894
rect 519502 452658 519586 452894
rect 519822 452658 553266 452894
rect 553502 452658 553586 452894
rect 553822 452658 587262 452894
rect 587498 452658 587582 452894
rect 587818 452658 592650 452894
rect -8726 452574 592650 452658
rect -8726 452338 -3894 452574
rect -3658 452338 -3574 452574
rect -3338 452338 9266 452574
rect 9502 452338 9586 452574
rect 9822 452338 43266 452574
rect 43502 452338 43586 452574
rect 43822 452338 77266 452574
rect 77502 452338 77586 452574
rect 77822 452338 111266 452574
rect 111502 452338 111586 452574
rect 111822 452338 145266 452574
rect 145502 452338 145586 452574
rect 145822 452338 179266 452574
rect 179502 452338 179586 452574
rect 179822 452338 213266 452574
rect 213502 452338 213586 452574
rect 213822 452338 247266 452574
rect 247502 452338 247586 452574
rect 247822 452338 281266 452574
rect 281502 452338 281586 452574
rect 281822 452338 315266 452574
rect 315502 452338 315586 452574
rect 315822 452338 349266 452574
rect 349502 452338 349586 452574
rect 349822 452338 383266 452574
rect 383502 452338 383586 452574
rect 383822 452338 417266 452574
rect 417502 452338 417586 452574
rect 417822 452338 451266 452574
rect 451502 452338 451586 452574
rect 451822 452338 485266 452574
rect 485502 452338 485586 452574
rect 485822 452338 519266 452574
rect 519502 452338 519586 452574
rect 519822 452338 553266 452574
rect 553502 452338 553586 452574
rect 553822 452338 587262 452574
rect 587498 452338 587582 452574
rect 587818 452338 592650 452574
rect -8726 452306 592650 452338
rect -8726 449174 592650 449206
rect -8726 448938 -2934 449174
rect -2698 448938 -2614 449174
rect -2378 448938 5546 449174
rect 5782 448938 5866 449174
rect 6102 448938 39546 449174
rect 39782 448938 39866 449174
rect 40102 448938 73546 449174
rect 73782 448938 73866 449174
rect 74102 448938 107546 449174
rect 107782 448938 107866 449174
rect 108102 448938 141546 449174
rect 141782 448938 141866 449174
rect 142102 448938 175546 449174
rect 175782 448938 175866 449174
rect 176102 448938 209546 449174
rect 209782 448938 209866 449174
rect 210102 448938 243546 449174
rect 243782 448938 243866 449174
rect 244102 448938 277546 449174
rect 277782 448938 277866 449174
rect 278102 448938 311546 449174
rect 311782 448938 311866 449174
rect 312102 448938 345546 449174
rect 345782 448938 345866 449174
rect 346102 448938 379546 449174
rect 379782 448938 379866 449174
rect 380102 448938 413546 449174
rect 413782 448938 413866 449174
rect 414102 448938 447546 449174
rect 447782 448938 447866 449174
rect 448102 448938 481546 449174
rect 481782 448938 481866 449174
rect 482102 448938 515546 449174
rect 515782 448938 515866 449174
rect 516102 448938 549546 449174
rect 549782 448938 549866 449174
rect 550102 448938 586302 449174
rect 586538 448938 586622 449174
rect 586858 448938 592650 449174
rect -8726 448854 592650 448938
rect -8726 448618 -2934 448854
rect -2698 448618 -2614 448854
rect -2378 448618 5546 448854
rect 5782 448618 5866 448854
rect 6102 448618 39546 448854
rect 39782 448618 39866 448854
rect 40102 448618 73546 448854
rect 73782 448618 73866 448854
rect 74102 448618 107546 448854
rect 107782 448618 107866 448854
rect 108102 448618 141546 448854
rect 141782 448618 141866 448854
rect 142102 448618 175546 448854
rect 175782 448618 175866 448854
rect 176102 448618 209546 448854
rect 209782 448618 209866 448854
rect 210102 448618 243546 448854
rect 243782 448618 243866 448854
rect 244102 448618 277546 448854
rect 277782 448618 277866 448854
rect 278102 448618 311546 448854
rect 311782 448618 311866 448854
rect 312102 448618 345546 448854
rect 345782 448618 345866 448854
rect 346102 448618 379546 448854
rect 379782 448618 379866 448854
rect 380102 448618 413546 448854
rect 413782 448618 413866 448854
rect 414102 448618 447546 448854
rect 447782 448618 447866 448854
rect 448102 448618 481546 448854
rect 481782 448618 481866 448854
rect 482102 448618 515546 448854
rect 515782 448618 515866 448854
rect 516102 448618 549546 448854
rect 549782 448618 549866 448854
rect 550102 448618 586302 448854
rect 586538 448618 586622 448854
rect 586858 448618 592650 448854
rect -8726 448586 592650 448618
rect -8726 445454 592650 445486
rect -8726 445218 -1974 445454
rect -1738 445218 -1654 445454
rect -1418 445218 1826 445454
rect 2062 445218 2146 445454
rect 2382 445218 35826 445454
rect 36062 445218 36146 445454
rect 36382 445218 69826 445454
rect 70062 445218 70146 445454
rect 70382 445218 103826 445454
rect 104062 445218 104146 445454
rect 104382 445218 137826 445454
rect 138062 445218 138146 445454
rect 138382 445218 171826 445454
rect 172062 445218 172146 445454
rect 172382 445218 205826 445454
rect 206062 445218 206146 445454
rect 206382 445218 239826 445454
rect 240062 445218 240146 445454
rect 240382 445218 273826 445454
rect 274062 445218 274146 445454
rect 274382 445218 307826 445454
rect 308062 445218 308146 445454
rect 308382 445218 341826 445454
rect 342062 445218 342146 445454
rect 342382 445218 375826 445454
rect 376062 445218 376146 445454
rect 376382 445218 409826 445454
rect 410062 445218 410146 445454
rect 410382 445218 443826 445454
rect 444062 445218 444146 445454
rect 444382 445218 477826 445454
rect 478062 445218 478146 445454
rect 478382 445218 511826 445454
rect 512062 445218 512146 445454
rect 512382 445218 545826 445454
rect 546062 445218 546146 445454
rect 546382 445218 579826 445454
rect 580062 445218 580146 445454
rect 580382 445218 585342 445454
rect 585578 445218 585662 445454
rect 585898 445218 592650 445454
rect -8726 445134 592650 445218
rect -8726 444898 -1974 445134
rect -1738 444898 -1654 445134
rect -1418 444898 1826 445134
rect 2062 444898 2146 445134
rect 2382 444898 35826 445134
rect 36062 444898 36146 445134
rect 36382 444898 69826 445134
rect 70062 444898 70146 445134
rect 70382 444898 103826 445134
rect 104062 444898 104146 445134
rect 104382 444898 137826 445134
rect 138062 444898 138146 445134
rect 138382 444898 171826 445134
rect 172062 444898 172146 445134
rect 172382 444898 205826 445134
rect 206062 444898 206146 445134
rect 206382 444898 239826 445134
rect 240062 444898 240146 445134
rect 240382 444898 273826 445134
rect 274062 444898 274146 445134
rect 274382 444898 307826 445134
rect 308062 444898 308146 445134
rect 308382 444898 341826 445134
rect 342062 444898 342146 445134
rect 342382 444898 375826 445134
rect 376062 444898 376146 445134
rect 376382 444898 409826 445134
rect 410062 444898 410146 445134
rect 410382 444898 443826 445134
rect 444062 444898 444146 445134
rect 444382 444898 477826 445134
rect 478062 444898 478146 445134
rect 478382 444898 511826 445134
rect 512062 444898 512146 445134
rect 512382 444898 545826 445134
rect 546062 444898 546146 445134
rect 546382 444898 579826 445134
rect 580062 444898 580146 445134
rect 580382 444898 585342 445134
rect 585578 444898 585662 445134
rect 585898 444898 592650 445134
rect -8726 444866 592650 444898
rect -8726 437494 592650 437526
rect -8726 437258 -8694 437494
rect -8458 437258 -8374 437494
rect -8138 437258 27866 437494
rect 28102 437258 28186 437494
rect 28422 437258 61866 437494
rect 62102 437258 62186 437494
rect 62422 437258 95866 437494
rect 96102 437258 96186 437494
rect 96422 437258 129866 437494
rect 130102 437258 130186 437494
rect 130422 437258 163866 437494
rect 164102 437258 164186 437494
rect 164422 437258 197866 437494
rect 198102 437258 198186 437494
rect 198422 437258 231866 437494
rect 232102 437258 232186 437494
rect 232422 437258 265866 437494
rect 266102 437258 266186 437494
rect 266422 437258 299866 437494
rect 300102 437258 300186 437494
rect 300422 437258 333866 437494
rect 334102 437258 334186 437494
rect 334422 437258 367866 437494
rect 368102 437258 368186 437494
rect 368422 437258 401866 437494
rect 402102 437258 402186 437494
rect 402422 437258 435866 437494
rect 436102 437258 436186 437494
rect 436422 437258 469866 437494
rect 470102 437258 470186 437494
rect 470422 437258 503866 437494
rect 504102 437258 504186 437494
rect 504422 437258 537866 437494
rect 538102 437258 538186 437494
rect 538422 437258 571866 437494
rect 572102 437258 572186 437494
rect 572422 437258 592062 437494
rect 592298 437258 592382 437494
rect 592618 437258 592650 437494
rect -8726 437174 592650 437258
rect -8726 436938 -8694 437174
rect -8458 436938 -8374 437174
rect -8138 436938 27866 437174
rect 28102 436938 28186 437174
rect 28422 436938 61866 437174
rect 62102 436938 62186 437174
rect 62422 436938 95866 437174
rect 96102 436938 96186 437174
rect 96422 436938 129866 437174
rect 130102 436938 130186 437174
rect 130422 436938 163866 437174
rect 164102 436938 164186 437174
rect 164422 436938 197866 437174
rect 198102 436938 198186 437174
rect 198422 436938 231866 437174
rect 232102 436938 232186 437174
rect 232422 436938 265866 437174
rect 266102 436938 266186 437174
rect 266422 436938 299866 437174
rect 300102 436938 300186 437174
rect 300422 436938 333866 437174
rect 334102 436938 334186 437174
rect 334422 436938 367866 437174
rect 368102 436938 368186 437174
rect 368422 436938 401866 437174
rect 402102 436938 402186 437174
rect 402422 436938 435866 437174
rect 436102 436938 436186 437174
rect 436422 436938 469866 437174
rect 470102 436938 470186 437174
rect 470422 436938 503866 437174
rect 504102 436938 504186 437174
rect 504422 436938 537866 437174
rect 538102 436938 538186 437174
rect 538422 436938 571866 437174
rect 572102 436938 572186 437174
rect 572422 436938 592062 437174
rect 592298 436938 592382 437174
rect 592618 436938 592650 437174
rect -8726 436906 592650 436938
rect -8726 433774 592650 433806
rect -8726 433538 -7734 433774
rect -7498 433538 -7414 433774
rect -7178 433538 24146 433774
rect 24382 433538 24466 433774
rect 24702 433538 58146 433774
rect 58382 433538 58466 433774
rect 58702 433538 92146 433774
rect 92382 433538 92466 433774
rect 92702 433538 126146 433774
rect 126382 433538 126466 433774
rect 126702 433538 160146 433774
rect 160382 433538 160466 433774
rect 160702 433538 194146 433774
rect 194382 433538 194466 433774
rect 194702 433538 228146 433774
rect 228382 433538 228466 433774
rect 228702 433538 262146 433774
rect 262382 433538 262466 433774
rect 262702 433538 296146 433774
rect 296382 433538 296466 433774
rect 296702 433538 330146 433774
rect 330382 433538 330466 433774
rect 330702 433538 364146 433774
rect 364382 433538 364466 433774
rect 364702 433538 398146 433774
rect 398382 433538 398466 433774
rect 398702 433538 432146 433774
rect 432382 433538 432466 433774
rect 432702 433538 466146 433774
rect 466382 433538 466466 433774
rect 466702 433538 500146 433774
rect 500382 433538 500466 433774
rect 500702 433538 534146 433774
rect 534382 433538 534466 433774
rect 534702 433538 568146 433774
rect 568382 433538 568466 433774
rect 568702 433538 591102 433774
rect 591338 433538 591422 433774
rect 591658 433538 592650 433774
rect -8726 433454 592650 433538
rect -8726 433218 -7734 433454
rect -7498 433218 -7414 433454
rect -7178 433218 24146 433454
rect 24382 433218 24466 433454
rect 24702 433218 58146 433454
rect 58382 433218 58466 433454
rect 58702 433218 92146 433454
rect 92382 433218 92466 433454
rect 92702 433218 126146 433454
rect 126382 433218 126466 433454
rect 126702 433218 160146 433454
rect 160382 433218 160466 433454
rect 160702 433218 194146 433454
rect 194382 433218 194466 433454
rect 194702 433218 228146 433454
rect 228382 433218 228466 433454
rect 228702 433218 262146 433454
rect 262382 433218 262466 433454
rect 262702 433218 296146 433454
rect 296382 433218 296466 433454
rect 296702 433218 330146 433454
rect 330382 433218 330466 433454
rect 330702 433218 364146 433454
rect 364382 433218 364466 433454
rect 364702 433218 398146 433454
rect 398382 433218 398466 433454
rect 398702 433218 432146 433454
rect 432382 433218 432466 433454
rect 432702 433218 466146 433454
rect 466382 433218 466466 433454
rect 466702 433218 500146 433454
rect 500382 433218 500466 433454
rect 500702 433218 534146 433454
rect 534382 433218 534466 433454
rect 534702 433218 568146 433454
rect 568382 433218 568466 433454
rect 568702 433218 591102 433454
rect 591338 433218 591422 433454
rect 591658 433218 592650 433454
rect -8726 433186 592650 433218
rect -8726 430054 592650 430086
rect -8726 429818 -6774 430054
rect -6538 429818 -6454 430054
rect -6218 429818 20426 430054
rect 20662 429818 20746 430054
rect 20982 429818 54426 430054
rect 54662 429818 54746 430054
rect 54982 429818 88426 430054
rect 88662 429818 88746 430054
rect 88982 429818 122426 430054
rect 122662 429818 122746 430054
rect 122982 429818 156426 430054
rect 156662 429818 156746 430054
rect 156982 429818 190426 430054
rect 190662 429818 190746 430054
rect 190982 429818 224426 430054
rect 224662 429818 224746 430054
rect 224982 429818 258426 430054
rect 258662 429818 258746 430054
rect 258982 429818 292426 430054
rect 292662 429818 292746 430054
rect 292982 429818 326426 430054
rect 326662 429818 326746 430054
rect 326982 429818 360426 430054
rect 360662 429818 360746 430054
rect 360982 429818 394426 430054
rect 394662 429818 394746 430054
rect 394982 429818 428426 430054
rect 428662 429818 428746 430054
rect 428982 429818 462426 430054
rect 462662 429818 462746 430054
rect 462982 429818 496426 430054
rect 496662 429818 496746 430054
rect 496982 429818 530426 430054
rect 530662 429818 530746 430054
rect 530982 429818 564426 430054
rect 564662 429818 564746 430054
rect 564982 429818 590142 430054
rect 590378 429818 590462 430054
rect 590698 429818 592650 430054
rect -8726 429734 592650 429818
rect -8726 429498 -6774 429734
rect -6538 429498 -6454 429734
rect -6218 429498 20426 429734
rect 20662 429498 20746 429734
rect 20982 429498 54426 429734
rect 54662 429498 54746 429734
rect 54982 429498 88426 429734
rect 88662 429498 88746 429734
rect 88982 429498 122426 429734
rect 122662 429498 122746 429734
rect 122982 429498 156426 429734
rect 156662 429498 156746 429734
rect 156982 429498 190426 429734
rect 190662 429498 190746 429734
rect 190982 429498 224426 429734
rect 224662 429498 224746 429734
rect 224982 429498 258426 429734
rect 258662 429498 258746 429734
rect 258982 429498 292426 429734
rect 292662 429498 292746 429734
rect 292982 429498 326426 429734
rect 326662 429498 326746 429734
rect 326982 429498 360426 429734
rect 360662 429498 360746 429734
rect 360982 429498 394426 429734
rect 394662 429498 394746 429734
rect 394982 429498 428426 429734
rect 428662 429498 428746 429734
rect 428982 429498 462426 429734
rect 462662 429498 462746 429734
rect 462982 429498 496426 429734
rect 496662 429498 496746 429734
rect 496982 429498 530426 429734
rect 530662 429498 530746 429734
rect 530982 429498 564426 429734
rect 564662 429498 564746 429734
rect 564982 429498 590142 429734
rect 590378 429498 590462 429734
rect 590698 429498 592650 429734
rect -8726 429466 592650 429498
rect -8726 426334 592650 426366
rect -8726 426098 -5814 426334
rect -5578 426098 -5494 426334
rect -5258 426098 16706 426334
rect 16942 426098 17026 426334
rect 17262 426098 50706 426334
rect 50942 426098 51026 426334
rect 51262 426098 84706 426334
rect 84942 426098 85026 426334
rect 85262 426098 118706 426334
rect 118942 426098 119026 426334
rect 119262 426098 152706 426334
rect 152942 426098 153026 426334
rect 153262 426098 186706 426334
rect 186942 426098 187026 426334
rect 187262 426098 220706 426334
rect 220942 426098 221026 426334
rect 221262 426098 254706 426334
rect 254942 426098 255026 426334
rect 255262 426098 288706 426334
rect 288942 426098 289026 426334
rect 289262 426098 322706 426334
rect 322942 426098 323026 426334
rect 323262 426098 356706 426334
rect 356942 426098 357026 426334
rect 357262 426098 390706 426334
rect 390942 426098 391026 426334
rect 391262 426098 424706 426334
rect 424942 426098 425026 426334
rect 425262 426098 458706 426334
rect 458942 426098 459026 426334
rect 459262 426098 492706 426334
rect 492942 426098 493026 426334
rect 493262 426098 526706 426334
rect 526942 426098 527026 426334
rect 527262 426098 560706 426334
rect 560942 426098 561026 426334
rect 561262 426098 589182 426334
rect 589418 426098 589502 426334
rect 589738 426098 592650 426334
rect -8726 426014 592650 426098
rect -8726 425778 -5814 426014
rect -5578 425778 -5494 426014
rect -5258 425778 16706 426014
rect 16942 425778 17026 426014
rect 17262 425778 50706 426014
rect 50942 425778 51026 426014
rect 51262 425778 84706 426014
rect 84942 425778 85026 426014
rect 85262 425778 118706 426014
rect 118942 425778 119026 426014
rect 119262 425778 152706 426014
rect 152942 425778 153026 426014
rect 153262 425778 186706 426014
rect 186942 425778 187026 426014
rect 187262 425778 220706 426014
rect 220942 425778 221026 426014
rect 221262 425778 254706 426014
rect 254942 425778 255026 426014
rect 255262 425778 288706 426014
rect 288942 425778 289026 426014
rect 289262 425778 322706 426014
rect 322942 425778 323026 426014
rect 323262 425778 356706 426014
rect 356942 425778 357026 426014
rect 357262 425778 390706 426014
rect 390942 425778 391026 426014
rect 391262 425778 424706 426014
rect 424942 425778 425026 426014
rect 425262 425778 458706 426014
rect 458942 425778 459026 426014
rect 459262 425778 492706 426014
rect 492942 425778 493026 426014
rect 493262 425778 526706 426014
rect 526942 425778 527026 426014
rect 527262 425778 560706 426014
rect 560942 425778 561026 426014
rect 561262 425778 589182 426014
rect 589418 425778 589502 426014
rect 589738 425778 592650 426014
rect -8726 425746 592650 425778
rect -8726 422614 592650 422646
rect -8726 422378 -4854 422614
rect -4618 422378 -4534 422614
rect -4298 422378 12986 422614
rect 13222 422378 13306 422614
rect 13542 422378 46986 422614
rect 47222 422378 47306 422614
rect 47542 422378 80986 422614
rect 81222 422378 81306 422614
rect 81542 422378 114986 422614
rect 115222 422378 115306 422614
rect 115542 422378 148986 422614
rect 149222 422378 149306 422614
rect 149542 422378 182986 422614
rect 183222 422378 183306 422614
rect 183542 422378 216986 422614
rect 217222 422378 217306 422614
rect 217542 422378 250986 422614
rect 251222 422378 251306 422614
rect 251542 422378 284986 422614
rect 285222 422378 285306 422614
rect 285542 422378 318986 422614
rect 319222 422378 319306 422614
rect 319542 422378 352986 422614
rect 353222 422378 353306 422614
rect 353542 422378 386986 422614
rect 387222 422378 387306 422614
rect 387542 422378 420986 422614
rect 421222 422378 421306 422614
rect 421542 422378 454986 422614
rect 455222 422378 455306 422614
rect 455542 422378 488986 422614
rect 489222 422378 489306 422614
rect 489542 422378 522986 422614
rect 523222 422378 523306 422614
rect 523542 422378 556986 422614
rect 557222 422378 557306 422614
rect 557542 422378 588222 422614
rect 588458 422378 588542 422614
rect 588778 422378 592650 422614
rect -8726 422294 592650 422378
rect -8726 422058 -4854 422294
rect -4618 422058 -4534 422294
rect -4298 422058 12986 422294
rect 13222 422058 13306 422294
rect 13542 422058 46986 422294
rect 47222 422058 47306 422294
rect 47542 422058 80986 422294
rect 81222 422058 81306 422294
rect 81542 422058 114986 422294
rect 115222 422058 115306 422294
rect 115542 422058 148986 422294
rect 149222 422058 149306 422294
rect 149542 422058 182986 422294
rect 183222 422058 183306 422294
rect 183542 422058 216986 422294
rect 217222 422058 217306 422294
rect 217542 422058 250986 422294
rect 251222 422058 251306 422294
rect 251542 422058 284986 422294
rect 285222 422058 285306 422294
rect 285542 422058 318986 422294
rect 319222 422058 319306 422294
rect 319542 422058 352986 422294
rect 353222 422058 353306 422294
rect 353542 422058 386986 422294
rect 387222 422058 387306 422294
rect 387542 422058 420986 422294
rect 421222 422058 421306 422294
rect 421542 422058 454986 422294
rect 455222 422058 455306 422294
rect 455542 422058 488986 422294
rect 489222 422058 489306 422294
rect 489542 422058 522986 422294
rect 523222 422058 523306 422294
rect 523542 422058 556986 422294
rect 557222 422058 557306 422294
rect 557542 422058 588222 422294
rect 588458 422058 588542 422294
rect 588778 422058 592650 422294
rect -8726 422026 592650 422058
rect -8726 418894 592650 418926
rect -8726 418658 -3894 418894
rect -3658 418658 -3574 418894
rect -3338 418658 9266 418894
rect 9502 418658 9586 418894
rect 9822 418658 43266 418894
rect 43502 418658 43586 418894
rect 43822 418658 77266 418894
rect 77502 418658 77586 418894
rect 77822 418658 111266 418894
rect 111502 418658 111586 418894
rect 111822 418658 145266 418894
rect 145502 418658 145586 418894
rect 145822 418658 179266 418894
rect 179502 418658 179586 418894
rect 179822 418658 213266 418894
rect 213502 418658 213586 418894
rect 213822 418658 247266 418894
rect 247502 418658 247586 418894
rect 247822 418658 281266 418894
rect 281502 418658 281586 418894
rect 281822 418658 315266 418894
rect 315502 418658 315586 418894
rect 315822 418658 349266 418894
rect 349502 418658 349586 418894
rect 349822 418658 383266 418894
rect 383502 418658 383586 418894
rect 383822 418658 417266 418894
rect 417502 418658 417586 418894
rect 417822 418658 451266 418894
rect 451502 418658 451586 418894
rect 451822 418658 485266 418894
rect 485502 418658 485586 418894
rect 485822 418658 519266 418894
rect 519502 418658 519586 418894
rect 519822 418658 553266 418894
rect 553502 418658 553586 418894
rect 553822 418658 587262 418894
rect 587498 418658 587582 418894
rect 587818 418658 592650 418894
rect -8726 418574 592650 418658
rect -8726 418338 -3894 418574
rect -3658 418338 -3574 418574
rect -3338 418338 9266 418574
rect 9502 418338 9586 418574
rect 9822 418338 43266 418574
rect 43502 418338 43586 418574
rect 43822 418338 77266 418574
rect 77502 418338 77586 418574
rect 77822 418338 111266 418574
rect 111502 418338 111586 418574
rect 111822 418338 145266 418574
rect 145502 418338 145586 418574
rect 145822 418338 179266 418574
rect 179502 418338 179586 418574
rect 179822 418338 213266 418574
rect 213502 418338 213586 418574
rect 213822 418338 247266 418574
rect 247502 418338 247586 418574
rect 247822 418338 281266 418574
rect 281502 418338 281586 418574
rect 281822 418338 315266 418574
rect 315502 418338 315586 418574
rect 315822 418338 349266 418574
rect 349502 418338 349586 418574
rect 349822 418338 383266 418574
rect 383502 418338 383586 418574
rect 383822 418338 417266 418574
rect 417502 418338 417586 418574
rect 417822 418338 451266 418574
rect 451502 418338 451586 418574
rect 451822 418338 485266 418574
rect 485502 418338 485586 418574
rect 485822 418338 519266 418574
rect 519502 418338 519586 418574
rect 519822 418338 553266 418574
rect 553502 418338 553586 418574
rect 553822 418338 587262 418574
rect 587498 418338 587582 418574
rect 587818 418338 592650 418574
rect -8726 418306 592650 418338
rect -8726 415174 592650 415206
rect -8726 414938 -2934 415174
rect -2698 414938 -2614 415174
rect -2378 414938 5546 415174
rect 5782 414938 5866 415174
rect 6102 414938 39546 415174
rect 39782 414938 39866 415174
rect 40102 414938 73546 415174
rect 73782 414938 73866 415174
rect 74102 414938 107546 415174
rect 107782 414938 107866 415174
rect 108102 414938 141546 415174
rect 141782 414938 141866 415174
rect 142102 414938 175546 415174
rect 175782 414938 175866 415174
rect 176102 414938 209546 415174
rect 209782 414938 209866 415174
rect 210102 414938 243546 415174
rect 243782 414938 243866 415174
rect 244102 414938 277546 415174
rect 277782 414938 277866 415174
rect 278102 414938 311546 415174
rect 311782 414938 311866 415174
rect 312102 414938 345546 415174
rect 345782 414938 345866 415174
rect 346102 414938 379546 415174
rect 379782 414938 379866 415174
rect 380102 414938 413546 415174
rect 413782 414938 413866 415174
rect 414102 414938 447546 415174
rect 447782 414938 447866 415174
rect 448102 414938 481546 415174
rect 481782 414938 481866 415174
rect 482102 414938 515546 415174
rect 515782 414938 515866 415174
rect 516102 414938 549546 415174
rect 549782 414938 549866 415174
rect 550102 414938 586302 415174
rect 586538 414938 586622 415174
rect 586858 414938 592650 415174
rect -8726 414854 592650 414938
rect -8726 414618 -2934 414854
rect -2698 414618 -2614 414854
rect -2378 414618 5546 414854
rect 5782 414618 5866 414854
rect 6102 414618 39546 414854
rect 39782 414618 39866 414854
rect 40102 414618 73546 414854
rect 73782 414618 73866 414854
rect 74102 414618 107546 414854
rect 107782 414618 107866 414854
rect 108102 414618 141546 414854
rect 141782 414618 141866 414854
rect 142102 414618 175546 414854
rect 175782 414618 175866 414854
rect 176102 414618 209546 414854
rect 209782 414618 209866 414854
rect 210102 414618 243546 414854
rect 243782 414618 243866 414854
rect 244102 414618 277546 414854
rect 277782 414618 277866 414854
rect 278102 414618 311546 414854
rect 311782 414618 311866 414854
rect 312102 414618 345546 414854
rect 345782 414618 345866 414854
rect 346102 414618 379546 414854
rect 379782 414618 379866 414854
rect 380102 414618 413546 414854
rect 413782 414618 413866 414854
rect 414102 414618 447546 414854
rect 447782 414618 447866 414854
rect 448102 414618 481546 414854
rect 481782 414618 481866 414854
rect 482102 414618 515546 414854
rect 515782 414618 515866 414854
rect 516102 414618 549546 414854
rect 549782 414618 549866 414854
rect 550102 414618 586302 414854
rect 586538 414618 586622 414854
rect 586858 414618 592650 414854
rect -8726 414586 592650 414618
rect -8726 411454 592650 411486
rect -8726 411218 -1974 411454
rect -1738 411218 -1654 411454
rect -1418 411218 1826 411454
rect 2062 411218 2146 411454
rect 2382 411218 35826 411454
rect 36062 411218 36146 411454
rect 36382 411218 69826 411454
rect 70062 411218 70146 411454
rect 70382 411218 103826 411454
rect 104062 411218 104146 411454
rect 104382 411218 137826 411454
rect 138062 411218 138146 411454
rect 138382 411218 171826 411454
rect 172062 411218 172146 411454
rect 172382 411218 205826 411454
rect 206062 411218 206146 411454
rect 206382 411218 239826 411454
rect 240062 411218 240146 411454
rect 240382 411218 273826 411454
rect 274062 411218 274146 411454
rect 274382 411218 307826 411454
rect 308062 411218 308146 411454
rect 308382 411218 341826 411454
rect 342062 411218 342146 411454
rect 342382 411218 375826 411454
rect 376062 411218 376146 411454
rect 376382 411218 409826 411454
rect 410062 411218 410146 411454
rect 410382 411218 443826 411454
rect 444062 411218 444146 411454
rect 444382 411218 477826 411454
rect 478062 411218 478146 411454
rect 478382 411218 511826 411454
rect 512062 411218 512146 411454
rect 512382 411218 545826 411454
rect 546062 411218 546146 411454
rect 546382 411218 579826 411454
rect 580062 411218 580146 411454
rect 580382 411218 585342 411454
rect 585578 411218 585662 411454
rect 585898 411218 592650 411454
rect -8726 411134 592650 411218
rect -8726 410898 -1974 411134
rect -1738 410898 -1654 411134
rect -1418 410898 1826 411134
rect 2062 410898 2146 411134
rect 2382 410898 35826 411134
rect 36062 410898 36146 411134
rect 36382 410898 69826 411134
rect 70062 410898 70146 411134
rect 70382 410898 103826 411134
rect 104062 410898 104146 411134
rect 104382 410898 137826 411134
rect 138062 410898 138146 411134
rect 138382 410898 171826 411134
rect 172062 410898 172146 411134
rect 172382 410898 205826 411134
rect 206062 410898 206146 411134
rect 206382 410898 239826 411134
rect 240062 410898 240146 411134
rect 240382 410898 273826 411134
rect 274062 410898 274146 411134
rect 274382 410898 307826 411134
rect 308062 410898 308146 411134
rect 308382 410898 341826 411134
rect 342062 410898 342146 411134
rect 342382 410898 375826 411134
rect 376062 410898 376146 411134
rect 376382 410898 409826 411134
rect 410062 410898 410146 411134
rect 410382 410898 443826 411134
rect 444062 410898 444146 411134
rect 444382 410898 477826 411134
rect 478062 410898 478146 411134
rect 478382 410898 511826 411134
rect 512062 410898 512146 411134
rect 512382 410898 545826 411134
rect 546062 410898 546146 411134
rect 546382 410898 579826 411134
rect 580062 410898 580146 411134
rect 580382 410898 585342 411134
rect 585578 410898 585662 411134
rect 585898 410898 592650 411134
rect -8726 410866 592650 410898
rect -8726 403494 592650 403526
rect -8726 403258 -8694 403494
rect -8458 403258 -8374 403494
rect -8138 403258 27866 403494
rect 28102 403258 28186 403494
rect 28422 403258 61866 403494
rect 62102 403258 62186 403494
rect 62422 403258 95866 403494
rect 96102 403258 96186 403494
rect 96422 403258 129866 403494
rect 130102 403258 130186 403494
rect 130422 403258 163866 403494
rect 164102 403258 164186 403494
rect 164422 403258 197866 403494
rect 198102 403258 198186 403494
rect 198422 403258 231866 403494
rect 232102 403258 232186 403494
rect 232422 403258 265866 403494
rect 266102 403258 266186 403494
rect 266422 403258 299866 403494
rect 300102 403258 300186 403494
rect 300422 403258 333866 403494
rect 334102 403258 334186 403494
rect 334422 403258 367866 403494
rect 368102 403258 368186 403494
rect 368422 403258 401866 403494
rect 402102 403258 402186 403494
rect 402422 403258 435866 403494
rect 436102 403258 436186 403494
rect 436422 403258 469866 403494
rect 470102 403258 470186 403494
rect 470422 403258 503866 403494
rect 504102 403258 504186 403494
rect 504422 403258 537866 403494
rect 538102 403258 538186 403494
rect 538422 403258 571866 403494
rect 572102 403258 572186 403494
rect 572422 403258 592062 403494
rect 592298 403258 592382 403494
rect 592618 403258 592650 403494
rect -8726 403174 592650 403258
rect -8726 402938 -8694 403174
rect -8458 402938 -8374 403174
rect -8138 402938 27866 403174
rect 28102 402938 28186 403174
rect 28422 402938 61866 403174
rect 62102 402938 62186 403174
rect 62422 402938 95866 403174
rect 96102 402938 96186 403174
rect 96422 402938 129866 403174
rect 130102 402938 130186 403174
rect 130422 402938 163866 403174
rect 164102 402938 164186 403174
rect 164422 402938 197866 403174
rect 198102 402938 198186 403174
rect 198422 402938 231866 403174
rect 232102 402938 232186 403174
rect 232422 402938 265866 403174
rect 266102 402938 266186 403174
rect 266422 402938 299866 403174
rect 300102 402938 300186 403174
rect 300422 402938 333866 403174
rect 334102 402938 334186 403174
rect 334422 402938 367866 403174
rect 368102 402938 368186 403174
rect 368422 402938 401866 403174
rect 402102 402938 402186 403174
rect 402422 402938 435866 403174
rect 436102 402938 436186 403174
rect 436422 402938 469866 403174
rect 470102 402938 470186 403174
rect 470422 402938 503866 403174
rect 504102 402938 504186 403174
rect 504422 402938 537866 403174
rect 538102 402938 538186 403174
rect 538422 402938 571866 403174
rect 572102 402938 572186 403174
rect 572422 402938 592062 403174
rect 592298 402938 592382 403174
rect 592618 402938 592650 403174
rect -8726 402906 592650 402938
rect -8726 399774 592650 399806
rect -8726 399538 -7734 399774
rect -7498 399538 -7414 399774
rect -7178 399538 24146 399774
rect 24382 399538 24466 399774
rect 24702 399538 58146 399774
rect 58382 399538 58466 399774
rect 58702 399538 92146 399774
rect 92382 399538 92466 399774
rect 92702 399538 126146 399774
rect 126382 399538 126466 399774
rect 126702 399538 160146 399774
rect 160382 399538 160466 399774
rect 160702 399538 194146 399774
rect 194382 399538 194466 399774
rect 194702 399538 228146 399774
rect 228382 399538 228466 399774
rect 228702 399538 262146 399774
rect 262382 399538 262466 399774
rect 262702 399538 296146 399774
rect 296382 399538 296466 399774
rect 296702 399538 330146 399774
rect 330382 399538 330466 399774
rect 330702 399538 364146 399774
rect 364382 399538 364466 399774
rect 364702 399538 398146 399774
rect 398382 399538 398466 399774
rect 398702 399538 432146 399774
rect 432382 399538 432466 399774
rect 432702 399538 466146 399774
rect 466382 399538 466466 399774
rect 466702 399538 500146 399774
rect 500382 399538 500466 399774
rect 500702 399538 534146 399774
rect 534382 399538 534466 399774
rect 534702 399538 568146 399774
rect 568382 399538 568466 399774
rect 568702 399538 591102 399774
rect 591338 399538 591422 399774
rect 591658 399538 592650 399774
rect -8726 399454 592650 399538
rect -8726 399218 -7734 399454
rect -7498 399218 -7414 399454
rect -7178 399218 24146 399454
rect 24382 399218 24466 399454
rect 24702 399218 58146 399454
rect 58382 399218 58466 399454
rect 58702 399218 92146 399454
rect 92382 399218 92466 399454
rect 92702 399218 126146 399454
rect 126382 399218 126466 399454
rect 126702 399218 160146 399454
rect 160382 399218 160466 399454
rect 160702 399218 194146 399454
rect 194382 399218 194466 399454
rect 194702 399218 228146 399454
rect 228382 399218 228466 399454
rect 228702 399218 262146 399454
rect 262382 399218 262466 399454
rect 262702 399218 296146 399454
rect 296382 399218 296466 399454
rect 296702 399218 330146 399454
rect 330382 399218 330466 399454
rect 330702 399218 364146 399454
rect 364382 399218 364466 399454
rect 364702 399218 398146 399454
rect 398382 399218 398466 399454
rect 398702 399218 432146 399454
rect 432382 399218 432466 399454
rect 432702 399218 466146 399454
rect 466382 399218 466466 399454
rect 466702 399218 500146 399454
rect 500382 399218 500466 399454
rect 500702 399218 534146 399454
rect 534382 399218 534466 399454
rect 534702 399218 568146 399454
rect 568382 399218 568466 399454
rect 568702 399218 591102 399454
rect 591338 399218 591422 399454
rect 591658 399218 592650 399454
rect -8726 399186 592650 399218
rect -8726 396054 592650 396086
rect -8726 395818 -6774 396054
rect -6538 395818 -6454 396054
rect -6218 395818 20426 396054
rect 20662 395818 20746 396054
rect 20982 395818 54426 396054
rect 54662 395818 54746 396054
rect 54982 395818 88426 396054
rect 88662 395818 88746 396054
rect 88982 395818 122426 396054
rect 122662 395818 122746 396054
rect 122982 395818 156426 396054
rect 156662 395818 156746 396054
rect 156982 395818 190426 396054
rect 190662 395818 190746 396054
rect 190982 395818 224426 396054
rect 224662 395818 224746 396054
rect 224982 395818 258426 396054
rect 258662 395818 258746 396054
rect 258982 395818 292426 396054
rect 292662 395818 292746 396054
rect 292982 395818 326426 396054
rect 326662 395818 326746 396054
rect 326982 395818 360426 396054
rect 360662 395818 360746 396054
rect 360982 395818 394426 396054
rect 394662 395818 394746 396054
rect 394982 395818 428426 396054
rect 428662 395818 428746 396054
rect 428982 395818 462426 396054
rect 462662 395818 462746 396054
rect 462982 395818 496426 396054
rect 496662 395818 496746 396054
rect 496982 395818 530426 396054
rect 530662 395818 530746 396054
rect 530982 395818 564426 396054
rect 564662 395818 564746 396054
rect 564982 395818 590142 396054
rect 590378 395818 590462 396054
rect 590698 395818 592650 396054
rect -8726 395734 592650 395818
rect -8726 395498 -6774 395734
rect -6538 395498 -6454 395734
rect -6218 395498 20426 395734
rect 20662 395498 20746 395734
rect 20982 395498 54426 395734
rect 54662 395498 54746 395734
rect 54982 395498 88426 395734
rect 88662 395498 88746 395734
rect 88982 395498 122426 395734
rect 122662 395498 122746 395734
rect 122982 395498 156426 395734
rect 156662 395498 156746 395734
rect 156982 395498 190426 395734
rect 190662 395498 190746 395734
rect 190982 395498 224426 395734
rect 224662 395498 224746 395734
rect 224982 395498 258426 395734
rect 258662 395498 258746 395734
rect 258982 395498 292426 395734
rect 292662 395498 292746 395734
rect 292982 395498 326426 395734
rect 326662 395498 326746 395734
rect 326982 395498 360426 395734
rect 360662 395498 360746 395734
rect 360982 395498 394426 395734
rect 394662 395498 394746 395734
rect 394982 395498 428426 395734
rect 428662 395498 428746 395734
rect 428982 395498 462426 395734
rect 462662 395498 462746 395734
rect 462982 395498 496426 395734
rect 496662 395498 496746 395734
rect 496982 395498 530426 395734
rect 530662 395498 530746 395734
rect 530982 395498 564426 395734
rect 564662 395498 564746 395734
rect 564982 395498 590142 395734
rect 590378 395498 590462 395734
rect 590698 395498 592650 395734
rect -8726 395466 592650 395498
rect -8726 392334 592650 392366
rect -8726 392098 -5814 392334
rect -5578 392098 -5494 392334
rect -5258 392098 16706 392334
rect 16942 392098 17026 392334
rect 17262 392098 50706 392334
rect 50942 392098 51026 392334
rect 51262 392098 84706 392334
rect 84942 392098 85026 392334
rect 85262 392098 118706 392334
rect 118942 392098 119026 392334
rect 119262 392098 152706 392334
rect 152942 392098 153026 392334
rect 153262 392098 186706 392334
rect 186942 392098 187026 392334
rect 187262 392098 220706 392334
rect 220942 392098 221026 392334
rect 221262 392098 254706 392334
rect 254942 392098 255026 392334
rect 255262 392098 288706 392334
rect 288942 392098 289026 392334
rect 289262 392098 322706 392334
rect 322942 392098 323026 392334
rect 323262 392098 356706 392334
rect 356942 392098 357026 392334
rect 357262 392098 390706 392334
rect 390942 392098 391026 392334
rect 391262 392098 424706 392334
rect 424942 392098 425026 392334
rect 425262 392098 458706 392334
rect 458942 392098 459026 392334
rect 459262 392098 492706 392334
rect 492942 392098 493026 392334
rect 493262 392098 526706 392334
rect 526942 392098 527026 392334
rect 527262 392098 560706 392334
rect 560942 392098 561026 392334
rect 561262 392098 589182 392334
rect 589418 392098 589502 392334
rect 589738 392098 592650 392334
rect -8726 392014 592650 392098
rect -8726 391778 -5814 392014
rect -5578 391778 -5494 392014
rect -5258 391778 16706 392014
rect 16942 391778 17026 392014
rect 17262 391778 50706 392014
rect 50942 391778 51026 392014
rect 51262 391778 84706 392014
rect 84942 391778 85026 392014
rect 85262 391778 118706 392014
rect 118942 391778 119026 392014
rect 119262 391778 152706 392014
rect 152942 391778 153026 392014
rect 153262 391778 186706 392014
rect 186942 391778 187026 392014
rect 187262 391778 220706 392014
rect 220942 391778 221026 392014
rect 221262 391778 254706 392014
rect 254942 391778 255026 392014
rect 255262 391778 288706 392014
rect 288942 391778 289026 392014
rect 289262 391778 322706 392014
rect 322942 391778 323026 392014
rect 323262 391778 356706 392014
rect 356942 391778 357026 392014
rect 357262 391778 390706 392014
rect 390942 391778 391026 392014
rect 391262 391778 424706 392014
rect 424942 391778 425026 392014
rect 425262 391778 458706 392014
rect 458942 391778 459026 392014
rect 459262 391778 492706 392014
rect 492942 391778 493026 392014
rect 493262 391778 526706 392014
rect 526942 391778 527026 392014
rect 527262 391778 560706 392014
rect 560942 391778 561026 392014
rect 561262 391778 589182 392014
rect 589418 391778 589502 392014
rect 589738 391778 592650 392014
rect -8726 391746 592650 391778
rect -8726 388614 592650 388646
rect -8726 388378 -4854 388614
rect -4618 388378 -4534 388614
rect -4298 388378 12986 388614
rect 13222 388378 13306 388614
rect 13542 388378 46986 388614
rect 47222 388378 47306 388614
rect 47542 388378 80986 388614
rect 81222 388378 81306 388614
rect 81542 388378 114986 388614
rect 115222 388378 115306 388614
rect 115542 388378 148986 388614
rect 149222 388378 149306 388614
rect 149542 388378 182986 388614
rect 183222 388378 183306 388614
rect 183542 388378 216986 388614
rect 217222 388378 217306 388614
rect 217542 388378 250986 388614
rect 251222 388378 251306 388614
rect 251542 388378 284986 388614
rect 285222 388378 285306 388614
rect 285542 388378 318986 388614
rect 319222 388378 319306 388614
rect 319542 388378 352986 388614
rect 353222 388378 353306 388614
rect 353542 388378 386986 388614
rect 387222 388378 387306 388614
rect 387542 388378 420986 388614
rect 421222 388378 421306 388614
rect 421542 388378 454986 388614
rect 455222 388378 455306 388614
rect 455542 388378 488986 388614
rect 489222 388378 489306 388614
rect 489542 388378 522986 388614
rect 523222 388378 523306 388614
rect 523542 388378 556986 388614
rect 557222 388378 557306 388614
rect 557542 388378 588222 388614
rect 588458 388378 588542 388614
rect 588778 388378 592650 388614
rect -8726 388294 592650 388378
rect -8726 388058 -4854 388294
rect -4618 388058 -4534 388294
rect -4298 388058 12986 388294
rect 13222 388058 13306 388294
rect 13542 388058 46986 388294
rect 47222 388058 47306 388294
rect 47542 388058 80986 388294
rect 81222 388058 81306 388294
rect 81542 388058 114986 388294
rect 115222 388058 115306 388294
rect 115542 388058 148986 388294
rect 149222 388058 149306 388294
rect 149542 388058 182986 388294
rect 183222 388058 183306 388294
rect 183542 388058 216986 388294
rect 217222 388058 217306 388294
rect 217542 388058 250986 388294
rect 251222 388058 251306 388294
rect 251542 388058 284986 388294
rect 285222 388058 285306 388294
rect 285542 388058 318986 388294
rect 319222 388058 319306 388294
rect 319542 388058 352986 388294
rect 353222 388058 353306 388294
rect 353542 388058 386986 388294
rect 387222 388058 387306 388294
rect 387542 388058 420986 388294
rect 421222 388058 421306 388294
rect 421542 388058 454986 388294
rect 455222 388058 455306 388294
rect 455542 388058 488986 388294
rect 489222 388058 489306 388294
rect 489542 388058 522986 388294
rect 523222 388058 523306 388294
rect 523542 388058 556986 388294
rect 557222 388058 557306 388294
rect 557542 388058 588222 388294
rect 588458 388058 588542 388294
rect 588778 388058 592650 388294
rect -8726 388026 592650 388058
rect -8726 384894 592650 384926
rect -8726 384658 -3894 384894
rect -3658 384658 -3574 384894
rect -3338 384658 9266 384894
rect 9502 384658 9586 384894
rect 9822 384658 43266 384894
rect 43502 384658 43586 384894
rect 43822 384658 77266 384894
rect 77502 384658 77586 384894
rect 77822 384658 111266 384894
rect 111502 384658 111586 384894
rect 111822 384658 145266 384894
rect 145502 384658 145586 384894
rect 145822 384658 179266 384894
rect 179502 384658 179586 384894
rect 179822 384658 213266 384894
rect 213502 384658 213586 384894
rect 213822 384658 247266 384894
rect 247502 384658 247586 384894
rect 247822 384658 281266 384894
rect 281502 384658 281586 384894
rect 281822 384658 315266 384894
rect 315502 384658 315586 384894
rect 315822 384658 349266 384894
rect 349502 384658 349586 384894
rect 349822 384658 383266 384894
rect 383502 384658 383586 384894
rect 383822 384658 417266 384894
rect 417502 384658 417586 384894
rect 417822 384658 451266 384894
rect 451502 384658 451586 384894
rect 451822 384658 485266 384894
rect 485502 384658 485586 384894
rect 485822 384658 519266 384894
rect 519502 384658 519586 384894
rect 519822 384658 553266 384894
rect 553502 384658 553586 384894
rect 553822 384658 587262 384894
rect 587498 384658 587582 384894
rect 587818 384658 592650 384894
rect -8726 384574 592650 384658
rect -8726 384338 -3894 384574
rect -3658 384338 -3574 384574
rect -3338 384338 9266 384574
rect 9502 384338 9586 384574
rect 9822 384338 43266 384574
rect 43502 384338 43586 384574
rect 43822 384338 77266 384574
rect 77502 384338 77586 384574
rect 77822 384338 111266 384574
rect 111502 384338 111586 384574
rect 111822 384338 145266 384574
rect 145502 384338 145586 384574
rect 145822 384338 179266 384574
rect 179502 384338 179586 384574
rect 179822 384338 213266 384574
rect 213502 384338 213586 384574
rect 213822 384338 247266 384574
rect 247502 384338 247586 384574
rect 247822 384338 281266 384574
rect 281502 384338 281586 384574
rect 281822 384338 315266 384574
rect 315502 384338 315586 384574
rect 315822 384338 349266 384574
rect 349502 384338 349586 384574
rect 349822 384338 383266 384574
rect 383502 384338 383586 384574
rect 383822 384338 417266 384574
rect 417502 384338 417586 384574
rect 417822 384338 451266 384574
rect 451502 384338 451586 384574
rect 451822 384338 485266 384574
rect 485502 384338 485586 384574
rect 485822 384338 519266 384574
rect 519502 384338 519586 384574
rect 519822 384338 553266 384574
rect 553502 384338 553586 384574
rect 553822 384338 587262 384574
rect 587498 384338 587582 384574
rect 587818 384338 592650 384574
rect -8726 384306 592650 384338
rect -8726 381174 592650 381206
rect -8726 380938 -2934 381174
rect -2698 380938 -2614 381174
rect -2378 380938 5546 381174
rect 5782 380938 5866 381174
rect 6102 380938 39546 381174
rect 39782 380938 39866 381174
rect 40102 380938 73546 381174
rect 73782 380938 73866 381174
rect 74102 380938 107546 381174
rect 107782 380938 107866 381174
rect 108102 380938 141546 381174
rect 141782 380938 141866 381174
rect 142102 380938 175546 381174
rect 175782 380938 175866 381174
rect 176102 380938 209546 381174
rect 209782 380938 209866 381174
rect 210102 380938 243546 381174
rect 243782 380938 243866 381174
rect 244102 380938 277546 381174
rect 277782 380938 277866 381174
rect 278102 380938 311546 381174
rect 311782 380938 311866 381174
rect 312102 380938 345546 381174
rect 345782 380938 345866 381174
rect 346102 380938 379546 381174
rect 379782 380938 379866 381174
rect 380102 380938 413546 381174
rect 413782 380938 413866 381174
rect 414102 380938 447546 381174
rect 447782 380938 447866 381174
rect 448102 380938 481546 381174
rect 481782 380938 481866 381174
rect 482102 380938 515546 381174
rect 515782 380938 515866 381174
rect 516102 380938 549546 381174
rect 549782 380938 549866 381174
rect 550102 380938 586302 381174
rect 586538 380938 586622 381174
rect 586858 380938 592650 381174
rect -8726 380854 592650 380938
rect -8726 380618 -2934 380854
rect -2698 380618 -2614 380854
rect -2378 380618 5546 380854
rect 5782 380618 5866 380854
rect 6102 380618 39546 380854
rect 39782 380618 39866 380854
rect 40102 380618 73546 380854
rect 73782 380618 73866 380854
rect 74102 380618 107546 380854
rect 107782 380618 107866 380854
rect 108102 380618 141546 380854
rect 141782 380618 141866 380854
rect 142102 380618 175546 380854
rect 175782 380618 175866 380854
rect 176102 380618 209546 380854
rect 209782 380618 209866 380854
rect 210102 380618 243546 380854
rect 243782 380618 243866 380854
rect 244102 380618 277546 380854
rect 277782 380618 277866 380854
rect 278102 380618 311546 380854
rect 311782 380618 311866 380854
rect 312102 380618 345546 380854
rect 345782 380618 345866 380854
rect 346102 380618 379546 380854
rect 379782 380618 379866 380854
rect 380102 380618 413546 380854
rect 413782 380618 413866 380854
rect 414102 380618 447546 380854
rect 447782 380618 447866 380854
rect 448102 380618 481546 380854
rect 481782 380618 481866 380854
rect 482102 380618 515546 380854
rect 515782 380618 515866 380854
rect 516102 380618 549546 380854
rect 549782 380618 549866 380854
rect 550102 380618 586302 380854
rect 586538 380618 586622 380854
rect 586858 380618 592650 380854
rect -8726 380586 592650 380618
rect -8726 377454 592650 377486
rect -8726 377218 -1974 377454
rect -1738 377218 -1654 377454
rect -1418 377218 1826 377454
rect 2062 377218 2146 377454
rect 2382 377218 35826 377454
rect 36062 377218 36146 377454
rect 36382 377218 69826 377454
rect 70062 377218 70146 377454
rect 70382 377218 103826 377454
rect 104062 377218 104146 377454
rect 104382 377218 137826 377454
rect 138062 377218 138146 377454
rect 138382 377218 171826 377454
rect 172062 377218 172146 377454
rect 172382 377218 205826 377454
rect 206062 377218 206146 377454
rect 206382 377218 239826 377454
rect 240062 377218 240146 377454
rect 240382 377218 273826 377454
rect 274062 377218 274146 377454
rect 274382 377218 307826 377454
rect 308062 377218 308146 377454
rect 308382 377218 341826 377454
rect 342062 377218 342146 377454
rect 342382 377218 375826 377454
rect 376062 377218 376146 377454
rect 376382 377218 409826 377454
rect 410062 377218 410146 377454
rect 410382 377218 443826 377454
rect 444062 377218 444146 377454
rect 444382 377218 477826 377454
rect 478062 377218 478146 377454
rect 478382 377218 511826 377454
rect 512062 377218 512146 377454
rect 512382 377218 545826 377454
rect 546062 377218 546146 377454
rect 546382 377218 579826 377454
rect 580062 377218 580146 377454
rect 580382 377218 585342 377454
rect 585578 377218 585662 377454
rect 585898 377218 592650 377454
rect -8726 377134 592650 377218
rect -8726 376898 -1974 377134
rect -1738 376898 -1654 377134
rect -1418 376898 1826 377134
rect 2062 376898 2146 377134
rect 2382 376898 35826 377134
rect 36062 376898 36146 377134
rect 36382 376898 69826 377134
rect 70062 376898 70146 377134
rect 70382 376898 103826 377134
rect 104062 376898 104146 377134
rect 104382 376898 137826 377134
rect 138062 376898 138146 377134
rect 138382 376898 171826 377134
rect 172062 376898 172146 377134
rect 172382 376898 205826 377134
rect 206062 376898 206146 377134
rect 206382 376898 239826 377134
rect 240062 376898 240146 377134
rect 240382 376898 273826 377134
rect 274062 376898 274146 377134
rect 274382 376898 307826 377134
rect 308062 376898 308146 377134
rect 308382 376898 341826 377134
rect 342062 376898 342146 377134
rect 342382 376898 375826 377134
rect 376062 376898 376146 377134
rect 376382 376898 409826 377134
rect 410062 376898 410146 377134
rect 410382 376898 443826 377134
rect 444062 376898 444146 377134
rect 444382 376898 477826 377134
rect 478062 376898 478146 377134
rect 478382 376898 511826 377134
rect 512062 376898 512146 377134
rect 512382 376898 545826 377134
rect 546062 376898 546146 377134
rect 546382 376898 579826 377134
rect 580062 376898 580146 377134
rect 580382 376898 585342 377134
rect 585578 376898 585662 377134
rect 585898 376898 592650 377134
rect -8726 376866 592650 376898
rect -8726 369494 592650 369526
rect -8726 369258 -8694 369494
rect -8458 369258 -8374 369494
rect -8138 369258 27866 369494
rect 28102 369258 28186 369494
rect 28422 369258 61866 369494
rect 62102 369258 62186 369494
rect 62422 369258 95866 369494
rect 96102 369258 96186 369494
rect 96422 369258 129866 369494
rect 130102 369258 130186 369494
rect 130422 369258 163866 369494
rect 164102 369258 164186 369494
rect 164422 369258 197866 369494
rect 198102 369258 198186 369494
rect 198422 369258 231866 369494
rect 232102 369258 232186 369494
rect 232422 369258 265866 369494
rect 266102 369258 266186 369494
rect 266422 369258 299866 369494
rect 300102 369258 300186 369494
rect 300422 369258 333866 369494
rect 334102 369258 334186 369494
rect 334422 369258 367866 369494
rect 368102 369258 368186 369494
rect 368422 369258 401866 369494
rect 402102 369258 402186 369494
rect 402422 369258 435866 369494
rect 436102 369258 436186 369494
rect 436422 369258 469866 369494
rect 470102 369258 470186 369494
rect 470422 369258 503866 369494
rect 504102 369258 504186 369494
rect 504422 369258 537866 369494
rect 538102 369258 538186 369494
rect 538422 369258 571866 369494
rect 572102 369258 572186 369494
rect 572422 369258 592062 369494
rect 592298 369258 592382 369494
rect 592618 369258 592650 369494
rect -8726 369174 592650 369258
rect -8726 368938 -8694 369174
rect -8458 368938 -8374 369174
rect -8138 368938 27866 369174
rect 28102 368938 28186 369174
rect 28422 368938 61866 369174
rect 62102 368938 62186 369174
rect 62422 368938 95866 369174
rect 96102 368938 96186 369174
rect 96422 368938 129866 369174
rect 130102 368938 130186 369174
rect 130422 368938 163866 369174
rect 164102 368938 164186 369174
rect 164422 368938 197866 369174
rect 198102 368938 198186 369174
rect 198422 368938 231866 369174
rect 232102 368938 232186 369174
rect 232422 368938 265866 369174
rect 266102 368938 266186 369174
rect 266422 368938 299866 369174
rect 300102 368938 300186 369174
rect 300422 368938 333866 369174
rect 334102 368938 334186 369174
rect 334422 368938 367866 369174
rect 368102 368938 368186 369174
rect 368422 368938 401866 369174
rect 402102 368938 402186 369174
rect 402422 368938 435866 369174
rect 436102 368938 436186 369174
rect 436422 368938 469866 369174
rect 470102 368938 470186 369174
rect 470422 368938 503866 369174
rect 504102 368938 504186 369174
rect 504422 368938 537866 369174
rect 538102 368938 538186 369174
rect 538422 368938 571866 369174
rect 572102 368938 572186 369174
rect 572422 368938 592062 369174
rect 592298 368938 592382 369174
rect 592618 368938 592650 369174
rect -8726 368906 592650 368938
rect -8726 365774 592650 365806
rect -8726 365538 -7734 365774
rect -7498 365538 -7414 365774
rect -7178 365538 24146 365774
rect 24382 365538 24466 365774
rect 24702 365538 58146 365774
rect 58382 365538 58466 365774
rect 58702 365538 92146 365774
rect 92382 365538 92466 365774
rect 92702 365538 126146 365774
rect 126382 365538 126466 365774
rect 126702 365538 160146 365774
rect 160382 365538 160466 365774
rect 160702 365538 194146 365774
rect 194382 365538 194466 365774
rect 194702 365538 228146 365774
rect 228382 365538 228466 365774
rect 228702 365538 262146 365774
rect 262382 365538 262466 365774
rect 262702 365538 296146 365774
rect 296382 365538 296466 365774
rect 296702 365538 330146 365774
rect 330382 365538 330466 365774
rect 330702 365538 364146 365774
rect 364382 365538 364466 365774
rect 364702 365538 398146 365774
rect 398382 365538 398466 365774
rect 398702 365538 432146 365774
rect 432382 365538 432466 365774
rect 432702 365538 466146 365774
rect 466382 365538 466466 365774
rect 466702 365538 500146 365774
rect 500382 365538 500466 365774
rect 500702 365538 534146 365774
rect 534382 365538 534466 365774
rect 534702 365538 568146 365774
rect 568382 365538 568466 365774
rect 568702 365538 591102 365774
rect 591338 365538 591422 365774
rect 591658 365538 592650 365774
rect -8726 365454 592650 365538
rect -8726 365218 -7734 365454
rect -7498 365218 -7414 365454
rect -7178 365218 24146 365454
rect 24382 365218 24466 365454
rect 24702 365218 58146 365454
rect 58382 365218 58466 365454
rect 58702 365218 92146 365454
rect 92382 365218 92466 365454
rect 92702 365218 126146 365454
rect 126382 365218 126466 365454
rect 126702 365218 160146 365454
rect 160382 365218 160466 365454
rect 160702 365218 194146 365454
rect 194382 365218 194466 365454
rect 194702 365218 228146 365454
rect 228382 365218 228466 365454
rect 228702 365218 262146 365454
rect 262382 365218 262466 365454
rect 262702 365218 296146 365454
rect 296382 365218 296466 365454
rect 296702 365218 330146 365454
rect 330382 365218 330466 365454
rect 330702 365218 364146 365454
rect 364382 365218 364466 365454
rect 364702 365218 398146 365454
rect 398382 365218 398466 365454
rect 398702 365218 432146 365454
rect 432382 365218 432466 365454
rect 432702 365218 466146 365454
rect 466382 365218 466466 365454
rect 466702 365218 500146 365454
rect 500382 365218 500466 365454
rect 500702 365218 534146 365454
rect 534382 365218 534466 365454
rect 534702 365218 568146 365454
rect 568382 365218 568466 365454
rect 568702 365218 591102 365454
rect 591338 365218 591422 365454
rect 591658 365218 592650 365454
rect -8726 365186 592650 365218
rect -8726 362054 592650 362086
rect -8726 361818 -6774 362054
rect -6538 361818 -6454 362054
rect -6218 361818 20426 362054
rect 20662 361818 20746 362054
rect 20982 361818 54426 362054
rect 54662 361818 54746 362054
rect 54982 361818 88426 362054
rect 88662 361818 88746 362054
rect 88982 361818 122426 362054
rect 122662 361818 122746 362054
rect 122982 361818 156426 362054
rect 156662 361818 156746 362054
rect 156982 361818 190426 362054
rect 190662 361818 190746 362054
rect 190982 361818 224426 362054
rect 224662 361818 224746 362054
rect 224982 361818 258426 362054
rect 258662 361818 258746 362054
rect 258982 361818 292426 362054
rect 292662 361818 292746 362054
rect 292982 361818 326426 362054
rect 326662 361818 326746 362054
rect 326982 361818 360426 362054
rect 360662 361818 360746 362054
rect 360982 361818 394426 362054
rect 394662 361818 394746 362054
rect 394982 361818 428426 362054
rect 428662 361818 428746 362054
rect 428982 361818 462426 362054
rect 462662 361818 462746 362054
rect 462982 361818 496426 362054
rect 496662 361818 496746 362054
rect 496982 361818 530426 362054
rect 530662 361818 530746 362054
rect 530982 361818 564426 362054
rect 564662 361818 564746 362054
rect 564982 361818 590142 362054
rect 590378 361818 590462 362054
rect 590698 361818 592650 362054
rect -8726 361734 592650 361818
rect -8726 361498 -6774 361734
rect -6538 361498 -6454 361734
rect -6218 361498 20426 361734
rect 20662 361498 20746 361734
rect 20982 361498 54426 361734
rect 54662 361498 54746 361734
rect 54982 361498 88426 361734
rect 88662 361498 88746 361734
rect 88982 361498 122426 361734
rect 122662 361498 122746 361734
rect 122982 361498 156426 361734
rect 156662 361498 156746 361734
rect 156982 361498 190426 361734
rect 190662 361498 190746 361734
rect 190982 361498 224426 361734
rect 224662 361498 224746 361734
rect 224982 361498 258426 361734
rect 258662 361498 258746 361734
rect 258982 361498 292426 361734
rect 292662 361498 292746 361734
rect 292982 361498 326426 361734
rect 326662 361498 326746 361734
rect 326982 361498 360426 361734
rect 360662 361498 360746 361734
rect 360982 361498 394426 361734
rect 394662 361498 394746 361734
rect 394982 361498 428426 361734
rect 428662 361498 428746 361734
rect 428982 361498 462426 361734
rect 462662 361498 462746 361734
rect 462982 361498 496426 361734
rect 496662 361498 496746 361734
rect 496982 361498 530426 361734
rect 530662 361498 530746 361734
rect 530982 361498 564426 361734
rect 564662 361498 564746 361734
rect 564982 361498 590142 361734
rect 590378 361498 590462 361734
rect 590698 361498 592650 361734
rect -8726 361466 592650 361498
rect -8726 358334 592650 358366
rect -8726 358098 -5814 358334
rect -5578 358098 -5494 358334
rect -5258 358098 16706 358334
rect 16942 358098 17026 358334
rect 17262 358098 50706 358334
rect 50942 358098 51026 358334
rect 51262 358098 84706 358334
rect 84942 358098 85026 358334
rect 85262 358098 118706 358334
rect 118942 358098 119026 358334
rect 119262 358098 152706 358334
rect 152942 358098 153026 358334
rect 153262 358098 186706 358334
rect 186942 358098 187026 358334
rect 187262 358098 220706 358334
rect 220942 358098 221026 358334
rect 221262 358098 254706 358334
rect 254942 358098 255026 358334
rect 255262 358098 288706 358334
rect 288942 358098 289026 358334
rect 289262 358098 322706 358334
rect 322942 358098 323026 358334
rect 323262 358098 356706 358334
rect 356942 358098 357026 358334
rect 357262 358098 390706 358334
rect 390942 358098 391026 358334
rect 391262 358098 424706 358334
rect 424942 358098 425026 358334
rect 425262 358098 458706 358334
rect 458942 358098 459026 358334
rect 459262 358098 492706 358334
rect 492942 358098 493026 358334
rect 493262 358098 526706 358334
rect 526942 358098 527026 358334
rect 527262 358098 560706 358334
rect 560942 358098 561026 358334
rect 561262 358098 589182 358334
rect 589418 358098 589502 358334
rect 589738 358098 592650 358334
rect -8726 358014 592650 358098
rect -8726 357778 -5814 358014
rect -5578 357778 -5494 358014
rect -5258 357778 16706 358014
rect 16942 357778 17026 358014
rect 17262 357778 50706 358014
rect 50942 357778 51026 358014
rect 51262 357778 84706 358014
rect 84942 357778 85026 358014
rect 85262 357778 118706 358014
rect 118942 357778 119026 358014
rect 119262 357778 152706 358014
rect 152942 357778 153026 358014
rect 153262 357778 186706 358014
rect 186942 357778 187026 358014
rect 187262 357778 220706 358014
rect 220942 357778 221026 358014
rect 221262 357778 254706 358014
rect 254942 357778 255026 358014
rect 255262 357778 288706 358014
rect 288942 357778 289026 358014
rect 289262 357778 322706 358014
rect 322942 357778 323026 358014
rect 323262 357778 356706 358014
rect 356942 357778 357026 358014
rect 357262 357778 390706 358014
rect 390942 357778 391026 358014
rect 391262 357778 424706 358014
rect 424942 357778 425026 358014
rect 425262 357778 458706 358014
rect 458942 357778 459026 358014
rect 459262 357778 492706 358014
rect 492942 357778 493026 358014
rect 493262 357778 526706 358014
rect 526942 357778 527026 358014
rect 527262 357778 560706 358014
rect 560942 357778 561026 358014
rect 561262 357778 589182 358014
rect 589418 357778 589502 358014
rect 589738 357778 592650 358014
rect -8726 357746 592650 357778
rect -8726 354614 592650 354646
rect -8726 354378 -4854 354614
rect -4618 354378 -4534 354614
rect -4298 354378 12986 354614
rect 13222 354378 13306 354614
rect 13542 354378 46986 354614
rect 47222 354378 47306 354614
rect 47542 354378 80986 354614
rect 81222 354378 81306 354614
rect 81542 354378 114986 354614
rect 115222 354378 115306 354614
rect 115542 354378 148986 354614
rect 149222 354378 149306 354614
rect 149542 354378 182986 354614
rect 183222 354378 183306 354614
rect 183542 354378 216986 354614
rect 217222 354378 217306 354614
rect 217542 354378 250986 354614
rect 251222 354378 251306 354614
rect 251542 354378 284986 354614
rect 285222 354378 285306 354614
rect 285542 354378 318986 354614
rect 319222 354378 319306 354614
rect 319542 354378 352986 354614
rect 353222 354378 353306 354614
rect 353542 354378 386986 354614
rect 387222 354378 387306 354614
rect 387542 354378 420986 354614
rect 421222 354378 421306 354614
rect 421542 354378 454986 354614
rect 455222 354378 455306 354614
rect 455542 354378 488986 354614
rect 489222 354378 489306 354614
rect 489542 354378 522986 354614
rect 523222 354378 523306 354614
rect 523542 354378 556986 354614
rect 557222 354378 557306 354614
rect 557542 354378 588222 354614
rect 588458 354378 588542 354614
rect 588778 354378 592650 354614
rect -8726 354294 592650 354378
rect -8726 354058 -4854 354294
rect -4618 354058 -4534 354294
rect -4298 354058 12986 354294
rect 13222 354058 13306 354294
rect 13542 354058 46986 354294
rect 47222 354058 47306 354294
rect 47542 354058 80986 354294
rect 81222 354058 81306 354294
rect 81542 354058 114986 354294
rect 115222 354058 115306 354294
rect 115542 354058 148986 354294
rect 149222 354058 149306 354294
rect 149542 354058 182986 354294
rect 183222 354058 183306 354294
rect 183542 354058 216986 354294
rect 217222 354058 217306 354294
rect 217542 354058 250986 354294
rect 251222 354058 251306 354294
rect 251542 354058 284986 354294
rect 285222 354058 285306 354294
rect 285542 354058 318986 354294
rect 319222 354058 319306 354294
rect 319542 354058 352986 354294
rect 353222 354058 353306 354294
rect 353542 354058 386986 354294
rect 387222 354058 387306 354294
rect 387542 354058 420986 354294
rect 421222 354058 421306 354294
rect 421542 354058 454986 354294
rect 455222 354058 455306 354294
rect 455542 354058 488986 354294
rect 489222 354058 489306 354294
rect 489542 354058 522986 354294
rect 523222 354058 523306 354294
rect 523542 354058 556986 354294
rect 557222 354058 557306 354294
rect 557542 354058 588222 354294
rect 588458 354058 588542 354294
rect 588778 354058 592650 354294
rect -8726 354026 592650 354058
rect -8726 350894 592650 350926
rect -8726 350658 -3894 350894
rect -3658 350658 -3574 350894
rect -3338 350658 9266 350894
rect 9502 350658 9586 350894
rect 9822 350658 43266 350894
rect 43502 350658 43586 350894
rect 43822 350658 77266 350894
rect 77502 350658 77586 350894
rect 77822 350658 111266 350894
rect 111502 350658 111586 350894
rect 111822 350658 145266 350894
rect 145502 350658 145586 350894
rect 145822 350658 179266 350894
rect 179502 350658 179586 350894
rect 179822 350658 213266 350894
rect 213502 350658 213586 350894
rect 213822 350658 247266 350894
rect 247502 350658 247586 350894
rect 247822 350658 281266 350894
rect 281502 350658 281586 350894
rect 281822 350658 315266 350894
rect 315502 350658 315586 350894
rect 315822 350658 349266 350894
rect 349502 350658 349586 350894
rect 349822 350658 383266 350894
rect 383502 350658 383586 350894
rect 383822 350658 417266 350894
rect 417502 350658 417586 350894
rect 417822 350658 451266 350894
rect 451502 350658 451586 350894
rect 451822 350658 485266 350894
rect 485502 350658 485586 350894
rect 485822 350658 519266 350894
rect 519502 350658 519586 350894
rect 519822 350658 553266 350894
rect 553502 350658 553586 350894
rect 553822 350658 587262 350894
rect 587498 350658 587582 350894
rect 587818 350658 592650 350894
rect -8726 350574 592650 350658
rect -8726 350338 -3894 350574
rect -3658 350338 -3574 350574
rect -3338 350338 9266 350574
rect 9502 350338 9586 350574
rect 9822 350338 43266 350574
rect 43502 350338 43586 350574
rect 43822 350338 77266 350574
rect 77502 350338 77586 350574
rect 77822 350338 111266 350574
rect 111502 350338 111586 350574
rect 111822 350338 145266 350574
rect 145502 350338 145586 350574
rect 145822 350338 179266 350574
rect 179502 350338 179586 350574
rect 179822 350338 213266 350574
rect 213502 350338 213586 350574
rect 213822 350338 247266 350574
rect 247502 350338 247586 350574
rect 247822 350338 281266 350574
rect 281502 350338 281586 350574
rect 281822 350338 315266 350574
rect 315502 350338 315586 350574
rect 315822 350338 349266 350574
rect 349502 350338 349586 350574
rect 349822 350338 383266 350574
rect 383502 350338 383586 350574
rect 383822 350338 417266 350574
rect 417502 350338 417586 350574
rect 417822 350338 451266 350574
rect 451502 350338 451586 350574
rect 451822 350338 485266 350574
rect 485502 350338 485586 350574
rect 485822 350338 519266 350574
rect 519502 350338 519586 350574
rect 519822 350338 553266 350574
rect 553502 350338 553586 350574
rect 553822 350338 587262 350574
rect 587498 350338 587582 350574
rect 587818 350338 592650 350574
rect -8726 350306 592650 350338
rect -8726 347174 592650 347206
rect -8726 346938 -2934 347174
rect -2698 346938 -2614 347174
rect -2378 346938 5546 347174
rect 5782 346938 5866 347174
rect 6102 346938 39546 347174
rect 39782 346938 39866 347174
rect 40102 346938 73546 347174
rect 73782 346938 73866 347174
rect 74102 346938 107546 347174
rect 107782 346938 107866 347174
rect 108102 346938 141546 347174
rect 141782 346938 141866 347174
rect 142102 346938 175546 347174
rect 175782 346938 175866 347174
rect 176102 346938 209546 347174
rect 209782 346938 209866 347174
rect 210102 346938 243546 347174
rect 243782 346938 243866 347174
rect 244102 346938 277546 347174
rect 277782 346938 277866 347174
rect 278102 346938 311546 347174
rect 311782 346938 311866 347174
rect 312102 346938 345546 347174
rect 345782 346938 345866 347174
rect 346102 346938 379546 347174
rect 379782 346938 379866 347174
rect 380102 346938 413546 347174
rect 413782 346938 413866 347174
rect 414102 346938 447546 347174
rect 447782 346938 447866 347174
rect 448102 346938 481546 347174
rect 481782 346938 481866 347174
rect 482102 346938 515546 347174
rect 515782 346938 515866 347174
rect 516102 346938 549546 347174
rect 549782 346938 549866 347174
rect 550102 346938 586302 347174
rect 586538 346938 586622 347174
rect 586858 346938 592650 347174
rect -8726 346854 592650 346938
rect -8726 346618 -2934 346854
rect -2698 346618 -2614 346854
rect -2378 346618 5546 346854
rect 5782 346618 5866 346854
rect 6102 346618 39546 346854
rect 39782 346618 39866 346854
rect 40102 346618 73546 346854
rect 73782 346618 73866 346854
rect 74102 346618 107546 346854
rect 107782 346618 107866 346854
rect 108102 346618 141546 346854
rect 141782 346618 141866 346854
rect 142102 346618 175546 346854
rect 175782 346618 175866 346854
rect 176102 346618 209546 346854
rect 209782 346618 209866 346854
rect 210102 346618 243546 346854
rect 243782 346618 243866 346854
rect 244102 346618 277546 346854
rect 277782 346618 277866 346854
rect 278102 346618 311546 346854
rect 311782 346618 311866 346854
rect 312102 346618 345546 346854
rect 345782 346618 345866 346854
rect 346102 346618 379546 346854
rect 379782 346618 379866 346854
rect 380102 346618 413546 346854
rect 413782 346618 413866 346854
rect 414102 346618 447546 346854
rect 447782 346618 447866 346854
rect 448102 346618 481546 346854
rect 481782 346618 481866 346854
rect 482102 346618 515546 346854
rect 515782 346618 515866 346854
rect 516102 346618 549546 346854
rect 549782 346618 549866 346854
rect 550102 346618 586302 346854
rect 586538 346618 586622 346854
rect 586858 346618 592650 346854
rect -8726 346586 592650 346618
rect -8726 343454 592650 343486
rect -8726 343218 -1974 343454
rect -1738 343218 -1654 343454
rect -1418 343218 1826 343454
rect 2062 343218 2146 343454
rect 2382 343218 35826 343454
rect 36062 343218 36146 343454
rect 36382 343218 69826 343454
rect 70062 343218 70146 343454
rect 70382 343218 103826 343454
rect 104062 343218 104146 343454
rect 104382 343218 137826 343454
rect 138062 343218 138146 343454
rect 138382 343218 171826 343454
rect 172062 343218 172146 343454
rect 172382 343218 205826 343454
rect 206062 343218 206146 343454
rect 206382 343218 239826 343454
rect 240062 343218 240146 343454
rect 240382 343218 273826 343454
rect 274062 343218 274146 343454
rect 274382 343218 307826 343454
rect 308062 343218 308146 343454
rect 308382 343218 341826 343454
rect 342062 343218 342146 343454
rect 342382 343218 375826 343454
rect 376062 343218 376146 343454
rect 376382 343218 409826 343454
rect 410062 343218 410146 343454
rect 410382 343218 443826 343454
rect 444062 343218 444146 343454
rect 444382 343218 477826 343454
rect 478062 343218 478146 343454
rect 478382 343218 511826 343454
rect 512062 343218 512146 343454
rect 512382 343218 545826 343454
rect 546062 343218 546146 343454
rect 546382 343218 579826 343454
rect 580062 343218 580146 343454
rect 580382 343218 585342 343454
rect 585578 343218 585662 343454
rect 585898 343218 592650 343454
rect -8726 343134 592650 343218
rect -8726 342898 -1974 343134
rect -1738 342898 -1654 343134
rect -1418 342898 1826 343134
rect 2062 342898 2146 343134
rect 2382 342898 35826 343134
rect 36062 342898 36146 343134
rect 36382 342898 69826 343134
rect 70062 342898 70146 343134
rect 70382 342898 103826 343134
rect 104062 342898 104146 343134
rect 104382 342898 137826 343134
rect 138062 342898 138146 343134
rect 138382 342898 171826 343134
rect 172062 342898 172146 343134
rect 172382 342898 205826 343134
rect 206062 342898 206146 343134
rect 206382 342898 239826 343134
rect 240062 342898 240146 343134
rect 240382 342898 273826 343134
rect 274062 342898 274146 343134
rect 274382 342898 307826 343134
rect 308062 342898 308146 343134
rect 308382 342898 341826 343134
rect 342062 342898 342146 343134
rect 342382 342898 375826 343134
rect 376062 342898 376146 343134
rect 376382 342898 409826 343134
rect 410062 342898 410146 343134
rect 410382 342898 443826 343134
rect 444062 342898 444146 343134
rect 444382 342898 477826 343134
rect 478062 342898 478146 343134
rect 478382 342898 511826 343134
rect 512062 342898 512146 343134
rect 512382 342898 545826 343134
rect 546062 342898 546146 343134
rect 546382 342898 579826 343134
rect 580062 342898 580146 343134
rect 580382 342898 585342 343134
rect 585578 342898 585662 343134
rect 585898 342898 592650 343134
rect -8726 342866 592650 342898
rect -8726 335494 592650 335526
rect -8726 335258 -8694 335494
rect -8458 335258 -8374 335494
rect -8138 335258 27866 335494
rect 28102 335258 28186 335494
rect 28422 335258 61866 335494
rect 62102 335258 62186 335494
rect 62422 335258 95866 335494
rect 96102 335258 96186 335494
rect 96422 335258 129866 335494
rect 130102 335258 130186 335494
rect 130422 335258 163866 335494
rect 164102 335258 164186 335494
rect 164422 335258 197866 335494
rect 198102 335258 198186 335494
rect 198422 335258 231866 335494
rect 232102 335258 232186 335494
rect 232422 335258 265866 335494
rect 266102 335258 266186 335494
rect 266422 335258 299866 335494
rect 300102 335258 300186 335494
rect 300422 335258 333866 335494
rect 334102 335258 334186 335494
rect 334422 335258 367866 335494
rect 368102 335258 368186 335494
rect 368422 335258 401866 335494
rect 402102 335258 402186 335494
rect 402422 335258 435866 335494
rect 436102 335258 436186 335494
rect 436422 335258 469866 335494
rect 470102 335258 470186 335494
rect 470422 335258 503866 335494
rect 504102 335258 504186 335494
rect 504422 335258 537866 335494
rect 538102 335258 538186 335494
rect 538422 335258 571866 335494
rect 572102 335258 572186 335494
rect 572422 335258 592062 335494
rect 592298 335258 592382 335494
rect 592618 335258 592650 335494
rect -8726 335174 592650 335258
rect -8726 334938 -8694 335174
rect -8458 334938 -8374 335174
rect -8138 334938 27866 335174
rect 28102 334938 28186 335174
rect 28422 334938 61866 335174
rect 62102 334938 62186 335174
rect 62422 334938 95866 335174
rect 96102 334938 96186 335174
rect 96422 334938 129866 335174
rect 130102 334938 130186 335174
rect 130422 334938 163866 335174
rect 164102 334938 164186 335174
rect 164422 334938 197866 335174
rect 198102 334938 198186 335174
rect 198422 334938 231866 335174
rect 232102 334938 232186 335174
rect 232422 334938 265866 335174
rect 266102 334938 266186 335174
rect 266422 334938 299866 335174
rect 300102 334938 300186 335174
rect 300422 334938 333866 335174
rect 334102 334938 334186 335174
rect 334422 334938 367866 335174
rect 368102 334938 368186 335174
rect 368422 334938 401866 335174
rect 402102 334938 402186 335174
rect 402422 334938 435866 335174
rect 436102 334938 436186 335174
rect 436422 334938 469866 335174
rect 470102 334938 470186 335174
rect 470422 334938 503866 335174
rect 504102 334938 504186 335174
rect 504422 334938 537866 335174
rect 538102 334938 538186 335174
rect 538422 334938 571866 335174
rect 572102 334938 572186 335174
rect 572422 334938 592062 335174
rect 592298 334938 592382 335174
rect 592618 334938 592650 335174
rect -8726 334906 592650 334938
rect -8726 331774 592650 331806
rect -8726 331538 -7734 331774
rect -7498 331538 -7414 331774
rect -7178 331538 24146 331774
rect 24382 331538 24466 331774
rect 24702 331538 58146 331774
rect 58382 331538 58466 331774
rect 58702 331538 92146 331774
rect 92382 331538 92466 331774
rect 92702 331538 126146 331774
rect 126382 331538 126466 331774
rect 126702 331538 160146 331774
rect 160382 331538 160466 331774
rect 160702 331538 194146 331774
rect 194382 331538 194466 331774
rect 194702 331538 228146 331774
rect 228382 331538 228466 331774
rect 228702 331538 262146 331774
rect 262382 331538 262466 331774
rect 262702 331538 296146 331774
rect 296382 331538 296466 331774
rect 296702 331538 330146 331774
rect 330382 331538 330466 331774
rect 330702 331538 364146 331774
rect 364382 331538 364466 331774
rect 364702 331538 398146 331774
rect 398382 331538 398466 331774
rect 398702 331538 432146 331774
rect 432382 331538 432466 331774
rect 432702 331538 466146 331774
rect 466382 331538 466466 331774
rect 466702 331538 500146 331774
rect 500382 331538 500466 331774
rect 500702 331538 534146 331774
rect 534382 331538 534466 331774
rect 534702 331538 568146 331774
rect 568382 331538 568466 331774
rect 568702 331538 591102 331774
rect 591338 331538 591422 331774
rect 591658 331538 592650 331774
rect -8726 331454 592650 331538
rect -8726 331218 -7734 331454
rect -7498 331218 -7414 331454
rect -7178 331218 24146 331454
rect 24382 331218 24466 331454
rect 24702 331218 58146 331454
rect 58382 331218 58466 331454
rect 58702 331218 92146 331454
rect 92382 331218 92466 331454
rect 92702 331218 126146 331454
rect 126382 331218 126466 331454
rect 126702 331218 160146 331454
rect 160382 331218 160466 331454
rect 160702 331218 194146 331454
rect 194382 331218 194466 331454
rect 194702 331218 228146 331454
rect 228382 331218 228466 331454
rect 228702 331218 262146 331454
rect 262382 331218 262466 331454
rect 262702 331218 296146 331454
rect 296382 331218 296466 331454
rect 296702 331218 330146 331454
rect 330382 331218 330466 331454
rect 330702 331218 364146 331454
rect 364382 331218 364466 331454
rect 364702 331218 398146 331454
rect 398382 331218 398466 331454
rect 398702 331218 432146 331454
rect 432382 331218 432466 331454
rect 432702 331218 466146 331454
rect 466382 331218 466466 331454
rect 466702 331218 500146 331454
rect 500382 331218 500466 331454
rect 500702 331218 534146 331454
rect 534382 331218 534466 331454
rect 534702 331218 568146 331454
rect 568382 331218 568466 331454
rect 568702 331218 591102 331454
rect 591338 331218 591422 331454
rect 591658 331218 592650 331454
rect -8726 331186 592650 331218
rect -8726 328054 592650 328086
rect -8726 327818 -6774 328054
rect -6538 327818 -6454 328054
rect -6218 327818 20426 328054
rect 20662 327818 20746 328054
rect 20982 327818 54426 328054
rect 54662 327818 54746 328054
rect 54982 327818 88426 328054
rect 88662 327818 88746 328054
rect 88982 327818 122426 328054
rect 122662 327818 122746 328054
rect 122982 327818 156426 328054
rect 156662 327818 156746 328054
rect 156982 327818 190426 328054
rect 190662 327818 190746 328054
rect 190982 327818 224426 328054
rect 224662 327818 224746 328054
rect 224982 327818 258426 328054
rect 258662 327818 258746 328054
rect 258982 327818 292426 328054
rect 292662 327818 292746 328054
rect 292982 327818 326426 328054
rect 326662 327818 326746 328054
rect 326982 327818 360426 328054
rect 360662 327818 360746 328054
rect 360982 327818 394426 328054
rect 394662 327818 394746 328054
rect 394982 327818 428426 328054
rect 428662 327818 428746 328054
rect 428982 327818 462426 328054
rect 462662 327818 462746 328054
rect 462982 327818 496426 328054
rect 496662 327818 496746 328054
rect 496982 327818 530426 328054
rect 530662 327818 530746 328054
rect 530982 327818 564426 328054
rect 564662 327818 564746 328054
rect 564982 327818 590142 328054
rect 590378 327818 590462 328054
rect 590698 327818 592650 328054
rect -8726 327734 592650 327818
rect -8726 327498 -6774 327734
rect -6538 327498 -6454 327734
rect -6218 327498 20426 327734
rect 20662 327498 20746 327734
rect 20982 327498 54426 327734
rect 54662 327498 54746 327734
rect 54982 327498 88426 327734
rect 88662 327498 88746 327734
rect 88982 327498 122426 327734
rect 122662 327498 122746 327734
rect 122982 327498 156426 327734
rect 156662 327498 156746 327734
rect 156982 327498 190426 327734
rect 190662 327498 190746 327734
rect 190982 327498 224426 327734
rect 224662 327498 224746 327734
rect 224982 327498 258426 327734
rect 258662 327498 258746 327734
rect 258982 327498 292426 327734
rect 292662 327498 292746 327734
rect 292982 327498 326426 327734
rect 326662 327498 326746 327734
rect 326982 327498 360426 327734
rect 360662 327498 360746 327734
rect 360982 327498 394426 327734
rect 394662 327498 394746 327734
rect 394982 327498 428426 327734
rect 428662 327498 428746 327734
rect 428982 327498 462426 327734
rect 462662 327498 462746 327734
rect 462982 327498 496426 327734
rect 496662 327498 496746 327734
rect 496982 327498 530426 327734
rect 530662 327498 530746 327734
rect 530982 327498 564426 327734
rect 564662 327498 564746 327734
rect 564982 327498 590142 327734
rect 590378 327498 590462 327734
rect 590698 327498 592650 327734
rect -8726 327466 592650 327498
rect -8726 324334 592650 324366
rect -8726 324098 -5814 324334
rect -5578 324098 -5494 324334
rect -5258 324098 16706 324334
rect 16942 324098 17026 324334
rect 17262 324098 50706 324334
rect 50942 324098 51026 324334
rect 51262 324098 84706 324334
rect 84942 324098 85026 324334
rect 85262 324098 118706 324334
rect 118942 324098 119026 324334
rect 119262 324098 152706 324334
rect 152942 324098 153026 324334
rect 153262 324098 186706 324334
rect 186942 324098 187026 324334
rect 187262 324098 220706 324334
rect 220942 324098 221026 324334
rect 221262 324098 254706 324334
rect 254942 324098 255026 324334
rect 255262 324098 288706 324334
rect 288942 324098 289026 324334
rect 289262 324098 322706 324334
rect 322942 324098 323026 324334
rect 323262 324098 356706 324334
rect 356942 324098 357026 324334
rect 357262 324098 390706 324334
rect 390942 324098 391026 324334
rect 391262 324098 424706 324334
rect 424942 324098 425026 324334
rect 425262 324098 458706 324334
rect 458942 324098 459026 324334
rect 459262 324098 492706 324334
rect 492942 324098 493026 324334
rect 493262 324098 526706 324334
rect 526942 324098 527026 324334
rect 527262 324098 560706 324334
rect 560942 324098 561026 324334
rect 561262 324098 589182 324334
rect 589418 324098 589502 324334
rect 589738 324098 592650 324334
rect -8726 324014 592650 324098
rect -8726 323778 -5814 324014
rect -5578 323778 -5494 324014
rect -5258 323778 16706 324014
rect 16942 323778 17026 324014
rect 17262 323778 50706 324014
rect 50942 323778 51026 324014
rect 51262 323778 84706 324014
rect 84942 323778 85026 324014
rect 85262 323778 118706 324014
rect 118942 323778 119026 324014
rect 119262 323778 152706 324014
rect 152942 323778 153026 324014
rect 153262 323778 186706 324014
rect 186942 323778 187026 324014
rect 187262 323778 220706 324014
rect 220942 323778 221026 324014
rect 221262 323778 254706 324014
rect 254942 323778 255026 324014
rect 255262 323778 288706 324014
rect 288942 323778 289026 324014
rect 289262 323778 322706 324014
rect 322942 323778 323026 324014
rect 323262 323778 356706 324014
rect 356942 323778 357026 324014
rect 357262 323778 390706 324014
rect 390942 323778 391026 324014
rect 391262 323778 424706 324014
rect 424942 323778 425026 324014
rect 425262 323778 458706 324014
rect 458942 323778 459026 324014
rect 459262 323778 492706 324014
rect 492942 323778 493026 324014
rect 493262 323778 526706 324014
rect 526942 323778 527026 324014
rect 527262 323778 560706 324014
rect 560942 323778 561026 324014
rect 561262 323778 589182 324014
rect 589418 323778 589502 324014
rect 589738 323778 592650 324014
rect -8726 323746 592650 323778
rect -8726 320614 592650 320646
rect -8726 320378 -4854 320614
rect -4618 320378 -4534 320614
rect -4298 320378 12986 320614
rect 13222 320378 13306 320614
rect 13542 320378 46986 320614
rect 47222 320378 47306 320614
rect 47542 320378 80986 320614
rect 81222 320378 81306 320614
rect 81542 320378 114986 320614
rect 115222 320378 115306 320614
rect 115542 320378 148986 320614
rect 149222 320378 149306 320614
rect 149542 320378 182986 320614
rect 183222 320378 183306 320614
rect 183542 320378 216986 320614
rect 217222 320378 217306 320614
rect 217542 320378 250986 320614
rect 251222 320378 251306 320614
rect 251542 320378 284986 320614
rect 285222 320378 285306 320614
rect 285542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 352986 320614
rect 353222 320378 353306 320614
rect 353542 320378 386986 320614
rect 387222 320378 387306 320614
rect 387542 320378 420986 320614
rect 421222 320378 421306 320614
rect 421542 320378 454986 320614
rect 455222 320378 455306 320614
rect 455542 320378 488986 320614
rect 489222 320378 489306 320614
rect 489542 320378 522986 320614
rect 523222 320378 523306 320614
rect 523542 320378 556986 320614
rect 557222 320378 557306 320614
rect 557542 320378 588222 320614
rect 588458 320378 588542 320614
rect 588778 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -4854 320294
rect -4618 320058 -4534 320294
rect -4298 320058 12986 320294
rect 13222 320058 13306 320294
rect 13542 320058 46986 320294
rect 47222 320058 47306 320294
rect 47542 320058 80986 320294
rect 81222 320058 81306 320294
rect 81542 320058 114986 320294
rect 115222 320058 115306 320294
rect 115542 320058 148986 320294
rect 149222 320058 149306 320294
rect 149542 320058 182986 320294
rect 183222 320058 183306 320294
rect 183542 320058 216986 320294
rect 217222 320058 217306 320294
rect 217542 320058 250986 320294
rect 251222 320058 251306 320294
rect 251542 320058 284986 320294
rect 285222 320058 285306 320294
rect 285542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 352986 320294
rect 353222 320058 353306 320294
rect 353542 320058 386986 320294
rect 387222 320058 387306 320294
rect 387542 320058 420986 320294
rect 421222 320058 421306 320294
rect 421542 320058 454986 320294
rect 455222 320058 455306 320294
rect 455542 320058 488986 320294
rect 489222 320058 489306 320294
rect 489542 320058 522986 320294
rect 523222 320058 523306 320294
rect 523542 320058 556986 320294
rect 557222 320058 557306 320294
rect 557542 320058 588222 320294
rect 588458 320058 588542 320294
rect 588778 320058 592650 320294
rect -8726 320026 592650 320058
rect -8726 316894 592650 316926
rect -8726 316658 -3894 316894
rect -3658 316658 -3574 316894
rect -3338 316658 9266 316894
rect 9502 316658 9586 316894
rect 9822 316658 43266 316894
rect 43502 316658 43586 316894
rect 43822 316658 77266 316894
rect 77502 316658 77586 316894
rect 77822 316658 111266 316894
rect 111502 316658 111586 316894
rect 111822 316658 145266 316894
rect 145502 316658 145586 316894
rect 145822 316658 179266 316894
rect 179502 316658 179586 316894
rect 179822 316658 213266 316894
rect 213502 316658 213586 316894
rect 213822 316658 247266 316894
rect 247502 316658 247586 316894
rect 247822 316658 281266 316894
rect 281502 316658 281586 316894
rect 281822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 349266 316894
rect 349502 316658 349586 316894
rect 349822 316658 383266 316894
rect 383502 316658 383586 316894
rect 383822 316658 417266 316894
rect 417502 316658 417586 316894
rect 417822 316658 451266 316894
rect 451502 316658 451586 316894
rect 451822 316658 485266 316894
rect 485502 316658 485586 316894
rect 485822 316658 519266 316894
rect 519502 316658 519586 316894
rect 519822 316658 553266 316894
rect 553502 316658 553586 316894
rect 553822 316658 587262 316894
rect 587498 316658 587582 316894
rect 587818 316658 592650 316894
rect -8726 316574 592650 316658
rect -8726 316338 -3894 316574
rect -3658 316338 -3574 316574
rect -3338 316338 9266 316574
rect 9502 316338 9586 316574
rect 9822 316338 43266 316574
rect 43502 316338 43586 316574
rect 43822 316338 77266 316574
rect 77502 316338 77586 316574
rect 77822 316338 111266 316574
rect 111502 316338 111586 316574
rect 111822 316338 145266 316574
rect 145502 316338 145586 316574
rect 145822 316338 179266 316574
rect 179502 316338 179586 316574
rect 179822 316338 213266 316574
rect 213502 316338 213586 316574
rect 213822 316338 247266 316574
rect 247502 316338 247586 316574
rect 247822 316338 281266 316574
rect 281502 316338 281586 316574
rect 281822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 349266 316574
rect 349502 316338 349586 316574
rect 349822 316338 383266 316574
rect 383502 316338 383586 316574
rect 383822 316338 417266 316574
rect 417502 316338 417586 316574
rect 417822 316338 451266 316574
rect 451502 316338 451586 316574
rect 451822 316338 485266 316574
rect 485502 316338 485586 316574
rect 485822 316338 519266 316574
rect 519502 316338 519586 316574
rect 519822 316338 553266 316574
rect 553502 316338 553586 316574
rect 553822 316338 587262 316574
rect 587498 316338 587582 316574
rect 587818 316338 592650 316574
rect -8726 316306 592650 316338
rect -8726 313174 592650 313206
rect -8726 312938 -2934 313174
rect -2698 312938 -2614 313174
rect -2378 312938 5546 313174
rect 5782 312938 5866 313174
rect 6102 312938 39546 313174
rect 39782 312938 39866 313174
rect 40102 312938 73546 313174
rect 73782 312938 73866 313174
rect 74102 312938 107546 313174
rect 107782 312938 107866 313174
rect 108102 312938 141546 313174
rect 141782 312938 141866 313174
rect 142102 312938 175546 313174
rect 175782 312938 175866 313174
rect 176102 312938 209546 313174
rect 209782 312938 209866 313174
rect 210102 312938 243546 313174
rect 243782 312938 243866 313174
rect 244102 312938 277546 313174
rect 277782 312938 277866 313174
rect 278102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 345546 313174
rect 345782 312938 345866 313174
rect 346102 312938 379546 313174
rect 379782 312938 379866 313174
rect 380102 312938 413546 313174
rect 413782 312938 413866 313174
rect 414102 312938 447546 313174
rect 447782 312938 447866 313174
rect 448102 312938 481546 313174
rect 481782 312938 481866 313174
rect 482102 312938 515546 313174
rect 515782 312938 515866 313174
rect 516102 312938 549546 313174
rect 549782 312938 549866 313174
rect 550102 312938 586302 313174
rect 586538 312938 586622 313174
rect 586858 312938 592650 313174
rect -8726 312854 592650 312938
rect -8726 312618 -2934 312854
rect -2698 312618 -2614 312854
rect -2378 312618 5546 312854
rect 5782 312618 5866 312854
rect 6102 312618 39546 312854
rect 39782 312618 39866 312854
rect 40102 312618 73546 312854
rect 73782 312618 73866 312854
rect 74102 312618 107546 312854
rect 107782 312618 107866 312854
rect 108102 312618 141546 312854
rect 141782 312618 141866 312854
rect 142102 312618 175546 312854
rect 175782 312618 175866 312854
rect 176102 312618 209546 312854
rect 209782 312618 209866 312854
rect 210102 312618 243546 312854
rect 243782 312618 243866 312854
rect 244102 312618 277546 312854
rect 277782 312618 277866 312854
rect 278102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 345546 312854
rect 345782 312618 345866 312854
rect 346102 312618 379546 312854
rect 379782 312618 379866 312854
rect 380102 312618 413546 312854
rect 413782 312618 413866 312854
rect 414102 312618 447546 312854
rect 447782 312618 447866 312854
rect 448102 312618 481546 312854
rect 481782 312618 481866 312854
rect 482102 312618 515546 312854
rect 515782 312618 515866 312854
rect 516102 312618 549546 312854
rect 549782 312618 549866 312854
rect 550102 312618 586302 312854
rect 586538 312618 586622 312854
rect 586858 312618 592650 312854
rect -8726 312586 592650 312618
rect -8726 309454 592650 309486
rect -8726 309218 -1974 309454
rect -1738 309218 -1654 309454
rect -1418 309218 1826 309454
rect 2062 309218 2146 309454
rect 2382 309218 35826 309454
rect 36062 309218 36146 309454
rect 36382 309218 69826 309454
rect 70062 309218 70146 309454
rect 70382 309218 103826 309454
rect 104062 309218 104146 309454
rect 104382 309218 137826 309454
rect 138062 309218 138146 309454
rect 138382 309218 171826 309454
rect 172062 309218 172146 309454
rect 172382 309218 205826 309454
rect 206062 309218 206146 309454
rect 206382 309218 239826 309454
rect 240062 309218 240146 309454
rect 240382 309218 273826 309454
rect 274062 309218 274146 309454
rect 274382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 341826 309454
rect 342062 309218 342146 309454
rect 342382 309218 375826 309454
rect 376062 309218 376146 309454
rect 376382 309218 409826 309454
rect 410062 309218 410146 309454
rect 410382 309218 443826 309454
rect 444062 309218 444146 309454
rect 444382 309218 477826 309454
rect 478062 309218 478146 309454
rect 478382 309218 511826 309454
rect 512062 309218 512146 309454
rect 512382 309218 545826 309454
rect 546062 309218 546146 309454
rect 546382 309218 579826 309454
rect 580062 309218 580146 309454
rect 580382 309218 585342 309454
rect 585578 309218 585662 309454
rect 585898 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -1974 309134
rect -1738 308898 -1654 309134
rect -1418 308898 1826 309134
rect 2062 308898 2146 309134
rect 2382 308898 35826 309134
rect 36062 308898 36146 309134
rect 36382 308898 69826 309134
rect 70062 308898 70146 309134
rect 70382 308898 103826 309134
rect 104062 308898 104146 309134
rect 104382 308898 137826 309134
rect 138062 308898 138146 309134
rect 138382 308898 171826 309134
rect 172062 308898 172146 309134
rect 172382 308898 205826 309134
rect 206062 308898 206146 309134
rect 206382 308898 239826 309134
rect 240062 308898 240146 309134
rect 240382 308898 273826 309134
rect 274062 308898 274146 309134
rect 274382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 341826 309134
rect 342062 308898 342146 309134
rect 342382 308898 375826 309134
rect 376062 308898 376146 309134
rect 376382 308898 409826 309134
rect 410062 308898 410146 309134
rect 410382 308898 443826 309134
rect 444062 308898 444146 309134
rect 444382 308898 477826 309134
rect 478062 308898 478146 309134
rect 478382 308898 511826 309134
rect 512062 308898 512146 309134
rect 512382 308898 545826 309134
rect 546062 308898 546146 309134
rect 546382 308898 579826 309134
rect 580062 308898 580146 309134
rect 580382 308898 585342 309134
rect 585578 308898 585662 309134
rect 585898 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 301494 592650 301526
rect -8726 301258 -8694 301494
rect -8458 301258 -8374 301494
rect -8138 301258 27866 301494
rect 28102 301258 28186 301494
rect 28422 301258 61866 301494
rect 62102 301258 62186 301494
rect 62422 301258 95866 301494
rect 96102 301258 96186 301494
rect 96422 301258 129866 301494
rect 130102 301258 130186 301494
rect 130422 301258 163866 301494
rect 164102 301258 164186 301494
rect 164422 301258 197866 301494
rect 198102 301258 198186 301494
rect 198422 301258 231866 301494
rect 232102 301258 232186 301494
rect 232422 301258 265866 301494
rect 266102 301258 266186 301494
rect 266422 301258 299866 301494
rect 300102 301258 300186 301494
rect 300422 301258 333866 301494
rect 334102 301258 334186 301494
rect 334422 301258 367866 301494
rect 368102 301258 368186 301494
rect 368422 301258 401866 301494
rect 402102 301258 402186 301494
rect 402422 301258 435866 301494
rect 436102 301258 436186 301494
rect 436422 301258 469866 301494
rect 470102 301258 470186 301494
rect 470422 301258 503866 301494
rect 504102 301258 504186 301494
rect 504422 301258 537866 301494
rect 538102 301258 538186 301494
rect 538422 301258 571866 301494
rect 572102 301258 572186 301494
rect 572422 301258 592062 301494
rect 592298 301258 592382 301494
rect 592618 301258 592650 301494
rect -8726 301174 592650 301258
rect -8726 300938 -8694 301174
rect -8458 300938 -8374 301174
rect -8138 300938 27866 301174
rect 28102 300938 28186 301174
rect 28422 300938 61866 301174
rect 62102 300938 62186 301174
rect 62422 300938 95866 301174
rect 96102 300938 96186 301174
rect 96422 300938 129866 301174
rect 130102 300938 130186 301174
rect 130422 300938 163866 301174
rect 164102 300938 164186 301174
rect 164422 300938 197866 301174
rect 198102 300938 198186 301174
rect 198422 300938 231866 301174
rect 232102 300938 232186 301174
rect 232422 300938 265866 301174
rect 266102 300938 266186 301174
rect 266422 300938 299866 301174
rect 300102 300938 300186 301174
rect 300422 300938 333866 301174
rect 334102 300938 334186 301174
rect 334422 300938 367866 301174
rect 368102 300938 368186 301174
rect 368422 300938 401866 301174
rect 402102 300938 402186 301174
rect 402422 300938 435866 301174
rect 436102 300938 436186 301174
rect 436422 300938 469866 301174
rect 470102 300938 470186 301174
rect 470422 300938 503866 301174
rect 504102 300938 504186 301174
rect 504422 300938 537866 301174
rect 538102 300938 538186 301174
rect 538422 300938 571866 301174
rect 572102 300938 572186 301174
rect 572422 300938 592062 301174
rect 592298 300938 592382 301174
rect 592618 300938 592650 301174
rect -8726 300906 592650 300938
rect -8726 297774 592650 297806
rect -8726 297538 -7734 297774
rect -7498 297538 -7414 297774
rect -7178 297538 24146 297774
rect 24382 297538 24466 297774
rect 24702 297538 58146 297774
rect 58382 297538 58466 297774
rect 58702 297538 92146 297774
rect 92382 297538 92466 297774
rect 92702 297538 126146 297774
rect 126382 297538 126466 297774
rect 126702 297538 160146 297774
rect 160382 297538 160466 297774
rect 160702 297538 194146 297774
rect 194382 297538 194466 297774
rect 194702 297538 228146 297774
rect 228382 297538 228466 297774
rect 228702 297538 262146 297774
rect 262382 297538 262466 297774
rect 262702 297538 296146 297774
rect 296382 297538 296466 297774
rect 296702 297538 330146 297774
rect 330382 297538 330466 297774
rect 330702 297538 364146 297774
rect 364382 297538 364466 297774
rect 364702 297538 398146 297774
rect 398382 297538 398466 297774
rect 398702 297538 432146 297774
rect 432382 297538 432466 297774
rect 432702 297538 466146 297774
rect 466382 297538 466466 297774
rect 466702 297538 500146 297774
rect 500382 297538 500466 297774
rect 500702 297538 534146 297774
rect 534382 297538 534466 297774
rect 534702 297538 568146 297774
rect 568382 297538 568466 297774
rect 568702 297538 591102 297774
rect 591338 297538 591422 297774
rect 591658 297538 592650 297774
rect -8726 297454 592650 297538
rect -8726 297218 -7734 297454
rect -7498 297218 -7414 297454
rect -7178 297218 24146 297454
rect 24382 297218 24466 297454
rect 24702 297218 58146 297454
rect 58382 297218 58466 297454
rect 58702 297218 92146 297454
rect 92382 297218 92466 297454
rect 92702 297218 126146 297454
rect 126382 297218 126466 297454
rect 126702 297218 160146 297454
rect 160382 297218 160466 297454
rect 160702 297218 194146 297454
rect 194382 297218 194466 297454
rect 194702 297218 228146 297454
rect 228382 297218 228466 297454
rect 228702 297218 262146 297454
rect 262382 297218 262466 297454
rect 262702 297218 296146 297454
rect 296382 297218 296466 297454
rect 296702 297218 330146 297454
rect 330382 297218 330466 297454
rect 330702 297218 364146 297454
rect 364382 297218 364466 297454
rect 364702 297218 398146 297454
rect 398382 297218 398466 297454
rect 398702 297218 432146 297454
rect 432382 297218 432466 297454
rect 432702 297218 466146 297454
rect 466382 297218 466466 297454
rect 466702 297218 500146 297454
rect 500382 297218 500466 297454
rect 500702 297218 534146 297454
rect 534382 297218 534466 297454
rect 534702 297218 568146 297454
rect 568382 297218 568466 297454
rect 568702 297218 591102 297454
rect 591338 297218 591422 297454
rect 591658 297218 592650 297454
rect -8726 297186 592650 297218
rect -8726 294054 592650 294086
rect -8726 293818 -6774 294054
rect -6538 293818 -6454 294054
rect -6218 293818 20426 294054
rect 20662 293818 20746 294054
rect 20982 293818 54426 294054
rect 54662 293818 54746 294054
rect 54982 293818 88426 294054
rect 88662 293818 88746 294054
rect 88982 293818 122426 294054
rect 122662 293818 122746 294054
rect 122982 293818 156426 294054
rect 156662 293818 156746 294054
rect 156982 293818 190426 294054
rect 190662 293818 190746 294054
rect 190982 293818 224426 294054
rect 224662 293818 224746 294054
rect 224982 293818 258426 294054
rect 258662 293818 258746 294054
rect 258982 293818 292426 294054
rect 292662 293818 292746 294054
rect 292982 293818 326426 294054
rect 326662 293818 326746 294054
rect 326982 293818 360426 294054
rect 360662 293818 360746 294054
rect 360982 293818 394426 294054
rect 394662 293818 394746 294054
rect 394982 293818 428426 294054
rect 428662 293818 428746 294054
rect 428982 293818 462426 294054
rect 462662 293818 462746 294054
rect 462982 293818 496426 294054
rect 496662 293818 496746 294054
rect 496982 293818 530426 294054
rect 530662 293818 530746 294054
rect 530982 293818 564426 294054
rect 564662 293818 564746 294054
rect 564982 293818 590142 294054
rect 590378 293818 590462 294054
rect 590698 293818 592650 294054
rect -8726 293734 592650 293818
rect -8726 293498 -6774 293734
rect -6538 293498 -6454 293734
rect -6218 293498 20426 293734
rect 20662 293498 20746 293734
rect 20982 293498 54426 293734
rect 54662 293498 54746 293734
rect 54982 293498 88426 293734
rect 88662 293498 88746 293734
rect 88982 293498 122426 293734
rect 122662 293498 122746 293734
rect 122982 293498 156426 293734
rect 156662 293498 156746 293734
rect 156982 293498 190426 293734
rect 190662 293498 190746 293734
rect 190982 293498 224426 293734
rect 224662 293498 224746 293734
rect 224982 293498 258426 293734
rect 258662 293498 258746 293734
rect 258982 293498 292426 293734
rect 292662 293498 292746 293734
rect 292982 293498 326426 293734
rect 326662 293498 326746 293734
rect 326982 293498 360426 293734
rect 360662 293498 360746 293734
rect 360982 293498 394426 293734
rect 394662 293498 394746 293734
rect 394982 293498 428426 293734
rect 428662 293498 428746 293734
rect 428982 293498 462426 293734
rect 462662 293498 462746 293734
rect 462982 293498 496426 293734
rect 496662 293498 496746 293734
rect 496982 293498 530426 293734
rect 530662 293498 530746 293734
rect 530982 293498 564426 293734
rect 564662 293498 564746 293734
rect 564982 293498 590142 293734
rect 590378 293498 590462 293734
rect 590698 293498 592650 293734
rect -8726 293466 592650 293498
rect -8726 290334 592650 290366
rect -8726 290098 -5814 290334
rect -5578 290098 -5494 290334
rect -5258 290098 16706 290334
rect 16942 290098 17026 290334
rect 17262 290098 50706 290334
rect 50942 290098 51026 290334
rect 51262 290098 84706 290334
rect 84942 290098 85026 290334
rect 85262 290098 118706 290334
rect 118942 290098 119026 290334
rect 119262 290098 152706 290334
rect 152942 290098 153026 290334
rect 153262 290098 186706 290334
rect 186942 290098 187026 290334
rect 187262 290098 220706 290334
rect 220942 290098 221026 290334
rect 221262 290098 254706 290334
rect 254942 290098 255026 290334
rect 255262 290098 288706 290334
rect 288942 290098 289026 290334
rect 289262 290098 322706 290334
rect 322942 290098 323026 290334
rect 323262 290098 356706 290334
rect 356942 290098 357026 290334
rect 357262 290098 390706 290334
rect 390942 290098 391026 290334
rect 391262 290098 424706 290334
rect 424942 290098 425026 290334
rect 425262 290098 458706 290334
rect 458942 290098 459026 290334
rect 459262 290098 492706 290334
rect 492942 290098 493026 290334
rect 493262 290098 526706 290334
rect 526942 290098 527026 290334
rect 527262 290098 560706 290334
rect 560942 290098 561026 290334
rect 561262 290098 589182 290334
rect 589418 290098 589502 290334
rect 589738 290098 592650 290334
rect -8726 290014 592650 290098
rect -8726 289778 -5814 290014
rect -5578 289778 -5494 290014
rect -5258 289778 16706 290014
rect 16942 289778 17026 290014
rect 17262 289778 50706 290014
rect 50942 289778 51026 290014
rect 51262 289778 84706 290014
rect 84942 289778 85026 290014
rect 85262 289778 118706 290014
rect 118942 289778 119026 290014
rect 119262 289778 152706 290014
rect 152942 289778 153026 290014
rect 153262 289778 186706 290014
rect 186942 289778 187026 290014
rect 187262 289778 220706 290014
rect 220942 289778 221026 290014
rect 221262 289778 254706 290014
rect 254942 289778 255026 290014
rect 255262 289778 288706 290014
rect 288942 289778 289026 290014
rect 289262 289778 322706 290014
rect 322942 289778 323026 290014
rect 323262 289778 356706 290014
rect 356942 289778 357026 290014
rect 357262 289778 390706 290014
rect 390942 289778 391026 290014
rect 391262 289778 424706 290014
rect 424942 289778 425026 290014
rect 425262 289778 458706 290014
rect 458942 289778 459026 290014
rect 459262 289778 492706 290014
rect 492942 289778 493026 290014
rect 493262 289778 526706 290014
rect 526942 289778 527026 290014
rect 527262 289778 560706 290014
rect 560942 289778 561026 290014
rect 561262 289778 589182 290014
rect 589418 289778 589502 290014
rect 589738 289778 592650 290014
rect -8726 289746 592650 289778
rect -8726 286614 592650 286646
rect -8726 286378 -4854 286614
rect -4618 286378 -4534 286614
rect -4298 286378 12986 286614
rect 13222 286378 13306 286614
rect 13542 286378 46986 286614
rect 47222 286378 47306 286614
rect 47542 286378 80986 286614
rect 81222 286378 81306 286614
rect 81542 286378 114986 286614
rect 115222 286378 115306 286614
rect 115542 286378 148986 286614
rect 149222 286378 149306 286614
rect 149542 286378 182986 286614
rect 183222 286378 183306 286614
rect 183542 286378 216986 286614
rect 217222 286378 217306 286614
rect 217542 286378 250986 286614
rect 251222 286378 251306 286614
rect 251542 286378 284986 286614
rect 285222 286378 285306 286614
rect 285542 286378 318986 286614
rect 319222 286378 319306 286614
rect 319542 286378 352986 286614
rect 353222 286378 353306 286614
rect 353542 286378 386986 286614
rect 387222 286378 387306 286614
rect 387542 286378 420986 286614
rect 421222 286378 421306 286614
rect 421542 286378 454986 286614
rect 455222 286378 455306 286614
rect 455542 286378 488986 286614
rect 489222 286378 489306 286614
rect 489542 286378 522986 286614
rect 523222 286378 523306 286614
rect 523542 286378 556986 286614
rect 557222 286378 557306 286614
rect 557542 286378 588222 286614
rect 588458 286378 588542 286614
rect 588778 286378 592650 286614
rect -8726 286294 592650 286378
rect -8726 286058 -4854 286294
rect -4618 286058 -4534 286294
rect -4298 286058 12986 286294
rect 13222 286058 13306 286294
rect 13542 286058 46986 286294
rect 47222 286058 47306 286294
rect 47542 286058 80986 286294
rect 81222 286058 81306 286294
rect 81542 286058 114986 286294
rect 115222 286058 115306 286294
rect 115542 286058 148986 286294
rect 149222 286058 149306 286294
rect 149542 286058 182986 286294
rect 183222 286058 183306 286294
rect 183542 286058 216986 286294
rect 217222 286058 217306 286294
rect 217542 286058 250986 286294
rect 251222 286058 251306 286294
rect 251542 286058 284986 286294
rect 285222 286058 285306 286294
rect 285542 286058 318986 286294
rect 319222 286058 319306 286294
rect 319542 286058 352986 286294
rect 353222 286058 353306 286294
rect 353542 286058 386986 286294
rect 387222 286058 387306 286294
rect 387542 286058 420986 286294
rect 421222 286058 421306 286294
rect 421542 286058 454986 286294
rect 455222 286058 455306 286294
rect 455542 286058 488986 286294
rect 489222 286058 489306 286294
rect 489542 286058 522986 286294
rect 523222 286058 523306 286294
rect 523542 286058 556986 286294
rect 557222 286058 557306 286294
rect 557542 286058 588222 286294
rect 588458 286058 588542 286294
rect 588778 286058 592650 286294
rect -8726 286026 592650 286058
rect -8726 282894 592650 282926
rect -8726 282658 -3894 282894
rect -3658 282658 -3574 282894
rect -3338 282658 9266 282894
rect 9502 282658 9586 282894
rect 9822 282658 43266 282894
rect 43502 282658 43586 282894
rect 43822 282658 77266 282894
rect 77502 282658 77586 282894
rect 77822 282658 111266 282894
rect 111502 282658 111586 282894
rect 111822 282658 145266 282894
rect 145502 282658 145586 282894
rect 145822 282658 179266 282894
rect 179502 282658 179586 282894
rect 179822 282658 213266 282894
rect 213502 282658 213586 282894
rect 213822 282658 247266 282894
rect 247502 282658 247586 282894
rect 247822 282658 281266 282894
rect 281502 282658 281586 282894
rect 281822 282658 315266 282894
rect 315502 282658 315586 282894
rect 315822 282658 349266 282894
rect 349502 282658 349586 282894
rect 349822 282658 383266 282894
rect 383502 282658 383586 282894
rect 383822 282658 417266 282894
rect 417502 282658 417586 282894
rect 417822 282658 451266 282894
rect 451502 282658 451586 282894
rect 451822 282658 485266 282894
rect 485502 282658 485586 282894
rect 485822 282658 519266 282894
rect 519502 282658 519586 282894
rect 519822 282658 553266 282894
rect 553502 282658 553586 282894
rect 553822 282658 587262 282894
rect 587498 282658 587582 282894
rect 587818 282658 592650 282894
rect -8726 282574 592650 282658
rect -8726 282338 -3894 282574
rect -3658 282338 -3574 282574
rect -3338 282338 9266 282574
rect 9502 282338 9586 282574
rect 9822 282338 43266 282574
rect 43502 282338 43586 282574
rect 43822 282338 77266 282574
rect 77502 282338 77586 282574
rect 77822 282338 111266 282574
rect 111502 282338 111586 282574
rect 111822 282338 145266 282574
rect 145502 282338 145586 282574
rect 145822 282338 179266 282574
rect 179502 282338 179586 282574
rect 179822 282338 213266 282574
rect 213502 282338 213586 282574
rect 213822 282338 247266 282574
rect 247502 282338 247586 282574
rect 247822 282338 281266 282574
rect 281502 282338 281586 282574
rect 281822 282338 315266 282574
rect 315502 282338 315586 282574
rect 315822 282338 349266 282574
rect 349502 282338 349586 282574
rect 349822 282338 383266 282574
rect 383502 282338 383586 282574
rect 383822 282338 417266 282574
rect 417502 282338 417586 282574
rect 417822 282338 451266 282574
rect 451502 282338 451586 282574
rect 451822 282338 485266 282574
rect 485502 282338 485586 282574
rect 485822 282338 519266 282574
rect 519502 282338 519586 282574
rect 519822 282338 553266 282574
rect 553502 282338 553586 282574
rect 553822 282338 587262 282574
rect 587498 282338 587582 282574
rect 587818 282338 592650 282574
rect -8726 282306 592650 282338
rect -8726 279174 592650 279206
rect -8726 278938 -2934 279174
rect -2698 278938 -2614 279174
rect -2378 278938 5546 279174
rect 5782 278938 5866 279174
rect 6102 278938 39546 279174
rect 39782 278938 39866 279174
rect 40102 278938 73546 279174
rect 73782 278938 73866 279174
rect 74102 278938 107546 279174
rect 107782 278938 107866 279174
rect 108102 278938 141546 279174
rect 141782 278938 141866 279174
rect 142102 278938 175546 279174
rect 175782 278938 175866 279174
rect 176102 278938 209546 279174
rect 209782 278938 209866 279174
rect 210102 278938 243546 279174
rect 243782 278938 243866 279174
rect 244102 278938 277546 279174
rect 277782 278938 277866 279174
rect 278102 278938 311546 279174
rect 311782 278938 311866 279174
rect 312102 278938 345546 279174
rect 345782 278938 345866 279174
rect 346102 278938 379546 279174
rect 379782 278938 379866 279174
rect 380102 278938 413546 279174
rect 413782 278938 413866 279174
rect 414102 278938 447546 279174
rect 447782 278938 447866 279174
rect 448102 278938 481546 279174
rect 481782 278938 481866 279174
rect 482102 278938 515546 279174
rect 515782 278938 515866 279174
rect 516102 278938 549546 279174
rect 549782 278938 549866 279174
rect 550102 278938 586302 279174
rect 586538 278938 586622 279174
rect 586858 278938 592650 279174
rect -8726 278854 592650 278938
rect -8726 278618 -2934 278854
rect -2698 278618 -2614 278854
rect -2378 278618 5546 278854
rect 5782 278618 5866 278854
rect 6102 278618 39546 278854
rect 39782 278618 39866 278854
rect 40102 278618 73546 278854
rect 73782 278618 73866 278854
rect 74102 278618 107546 278854
rect 107782 278618 107866 278854
rect 108102 278618 141546 278854
rect 141782 278618 141866 278854
rect 142102 278618 175546 278854
rect 175782 278618 175866 278854
rect 176102 278618 209546 278854
rect 209782 278618 209866 278854
rect 210102 278618 243546 278854
rect 243782 278618 243866 278854
rect 244102 278618 277546 278854
rect 277782 278618 277866 278854
rect 278102 278618 311546 278854
rect 311782 278618 311866 278854
rect 312102 278618 345546 278854
rect 345782 278618 345866 278854
rect 346102 278618 379546 278854
rect 379782 278618 379866 278854
rect 380102 278618 413546 278854
rect 413782 278618 413866 278854
rect 414102 278618 447546 278854
rect 447782 278618 447866 278854
rect 448102 278618 481546 278854
rect 481782 278618 481866 278854
rect 482102 278618 515546 278854
rect 515782 278618 515866 278854
rect 516102 278618 549546 278854
rect 549782 278618 549866 278854
rect 550102 278618 586302 278854
rect 586538 278618 586622 278854
rect 586858 278618 592650 278854
rect -8726 278586 592650 278618
rect -8726 275454 592650 275486
rect -8726 275218 -1974 275454
rect -1738 275218 -1654 275454
rect -1418 275218 1826 275454
rect 2062 275218 2146 275454
rect 2382 275218 35826 275454
rect 36062 275218 36146 275454
rect 36382 275218 69826 275454
rect 70062 275218 70146 275454
rect 70382 275218 103826 275454
rect 104062 275218 104146 275454
rect 104382 275218 137826 275454
rect 138062 275218 138146 275454
rect 138382 275218 171826 275454
rect 172062 275218 172146 275454
rect 172382 275218 205826 275454
rect 206062 275218 206146 275454
rect 206382 275218 239826 275454
rect 240062 275218 240146 275454
rect 240382 275218 273826 275454
rect 274062 275218 274146 275454
rect 274382 275218 307826 275454
rect 308062 275218 308146 275454
rect 308382 275218 341826 275454
rect 342062 275218 342146 275454
rect 342382 275218 375826 275454
rect 376062 275218 376146 275454
rect 376382 275218 409826 275454
rect 410062 275218 410146 275454
rect 410382 275218 443826 275454
rect 444062 275218 444146 275454
rect 444382 275218 477826 275454
rect 478062 275218 478146 275454
rect 478382 275218 511826 275454
rect 512062 275218 512146 275454
rect 512382 275218 545826 275454
rect 546062 275218 546146 275454
rect 546382 275218 579826 275454
rect 580062 275218 580146 275454
rect 580382 275218 585342 275454
rect 585578 275218 585662 275454
rect 585898 275218 592650 275454
rect -8726 275134 592650 275218
rect -8726 274898 -1974 275134
rect -1738 274898 -1654 275134
rect -1418 274898 1826 275134
rect 2062 274898 2146 275134
rect 2382 274898 35826 275134
rect 36062 274898 36146 275134
rect 36382 274898 69826 275134
rect 70062 274898 70146 275134
rect 70382 274898 103826 275134
rect 104062 274898 104146 275134
rect 104382 274898 137826 275134
rect 138062 274898 138146 275134
rect 138382 274898 171826 275134
rect 172062 274898 172146 275134
rect 172382 274898 205826 275134
rect 206062 274898 206146 275134
rect 206382 274898 239826 275134
rect 240062 274898 240146 275134
rect 240382 274898 273826 275134
rect 274062 274898 274146 275134
rect 274382 274898 307826 275134
rect 308062 274898 308146 275134
rect 308382 274898 341826 275134
rect 342062 274898 342146 275134
rect 342382 274898 375826 275134
rect 376062 274898 376146 275134
rect 376382 274898 409826 275134
rect 410062 274898 410146 275134
rect 410382 274898 443826 275134
rect 444062 274898 444146 275134
rect 444382 274898 477826 275134
rect 478062 274898 478146 275134
rect 478382 274898 511826 275134
rect 512062 274898 512146 275134
rect 512382 274898 545826 275134
rect 546062 274898 546146 275134
rect 546382 274898 579826 275134
rect 580062 274898 580146 275134
rect 580382 274898 585342 275134
rect 585578 274898 585662 275134
rect 585898 274898 592650 275134
rect -8726 274866 592650 274898
rect -8726 267494 592650 267526
rect -8726 267258 -8694 267494
rect -8458 267258 -8374 267494
rect -8138 267258 27866 267494
rect 28102 267258 28186 267494
rect 28422 267258 61866 267494
rect 62102 267258 62186 267494
rect 62422 267258 95866 267494
rect 96102 267258 96186 267494
rect 96422 267258 129866 267494
rect 130102 267258 130186 267494
rect 130422 267258 163866 267494
rect 164102 267258 164186 267494
rect 164422 267258 197866 267494
rect 198102 267258 198186 267494
rect 198422 267258 231866 267494
rect 232102 267258 232186 267494
rect 232422 267258 265866 267494
rect 266102 267258 266186 267494
rect 266422 267258 299866 267494
rect 300102 267258 300186 267494
rect 300422 267258 333866 267494
rect 334102 267258 334186 267494
rect 334422 267258 367866 267494
rect 368102 267258 368186 267494
rect 368422 267258 401866 267494
rect 402102 267258 402186 267494
rect 402422 267258 435866 267494
rect 436102 267258 436186 267494
rect 436422 267258 469866 267494
rect 470102 267258 470186 267494
rect 470422 267258 503866 267494
rect 504102 267258 504186 267494
rect 504422 267258 537866 267494
rect 538102 267258 538186 267494
rect 538422 267258 571866 267494
rect 572102 267258 572186 267494
rect 572422 267258 592062 267494
rect 592298 267258 592382 267494
rect 592618 267258 592650 267494
rect -8726 267174 592650 267258
rect -8726 266938 -8694 267174
rect -8458 266938 -8374 267174
rect -8138 266938 27866 267174
rect 28102 266938 28186 267174
rect 28422 266938 61866 267174
rect 62102 266938 62186 267174
rect 62422 266938 95866 267174
rect 96102 266938 96186 267174
rect 96422 266938 129866 267174
rect 130102 266938 130186 267174
rect 130422 266938 163866 267174
rect 164102 266938 164186 267174
rect 164422 266938 197866 267174
rect 198102 266938 198186 267174
rect 198422 266938 231866 267174
rect 232102 266938 232186 267174
rect 232422 266938 265866 267174
rect 266102 266938 266186 267174
rect 266422 266938 299866 267174
rect 300102 266938 300186 267174
rect 300422 266938 333866 267174
rect 334102 266938 334186 267174
rect 334422 266938 367866 267174
rect 368102 266938 368186 267174
rect 368422 266938 401866 267174
rect 402102 266938 402186 267174
rect 402422 266938 435866 267174
rect 436102 266938 436186 267174
rect 436422 266938 469866 267174
rect 470102 266938 470186 267174
rect 470422 266938 503866 267174
rect 504102 266938 504186 267174
rect 504422 266938 537866 267174
rect 538102 266938 538186 267174
rect 538422 266938 571866 267174
rect 572102 266938 572186 267174
rect 572422 266938 592062 267174
rect 592298 266938 592382 267174
rect 592618 266938 592650 267174
rect -8726 266906 592650 266938
rect -8726 263774 592650 263806
rect -8726 263538 -7734 263774
rect -7498 263538 -7414 263774
rect -7178 263538 24146 263774
rect 24382 263538 24466 263774
rect 24702 263538 58146 263774
rect 58382 263538 58466 263774
rect 58702 263538 92146 263774
rect 92382 263538 92466 263774
rect 92702 263538 126146 263774
rect 126382 263538 126466 263774
rect 126702 263538 160146 263774
rect 160382 263538 160466 263774
rect 160702 263538 194146 263774
rect 194382 263538 194466 263774
rect 194702 263538 228146 263774
rect 228382 263538 228466 263774
rect 228702 263538 262146 263774
rect 262382 263538 262466 263774
rect 262702 263538 296146 263774
rect 296382 263538 296466 263774
rect 296702 263538 330146 263774
rect 330382 263538 330466 263774
rect 330702 263538 364146 263774
rect 364382 263538 364466 263774
rect 364702 263538 398146 263774
rect 398382 263538 398466 263774
rect 398702 263538 432146 263774
rect 432382 263538 432466 263774
rect 432702 263538 466146 263774
rect 466382 263538 466466 263774
rect 466702 263538 500146 263774
rect 500382 263538 500466 263774
rect 500702 263538 534146 263774
rect 534382 263538 534466 263774
rect 534702 263538 568146 263774
rect 568382 263538 568466 263774
rect 568702 263538 591102 263774
rect 591338 263538 591422 263774
rect 591658 263538 592650 263774
rect -8726 263454 592650 263538
rect -8726 263218 -7734 263454
rect -7498 263218 -7414 263454
rect -7178 263218 24146 263454
rect 24382 263218 24466 263454
rect 24702 263218 58146 263454
rect 58382 263218 58466 263454
rect 58702 263218 92146 263454
rect 92382 263218 92466 263454
rect 92702 263218 126146 263454
rect 126382 263218 126466 263454
rect 126702 263218 160146 263454
rect 160382 263218 160466 263454
rect 160702 263218 194146 263454
rect 194382 263218 194466 263454
rect 194702 263218 228146 263454
rect 228382 263218 228466 263454
rect 228702 263218 262146 263454
rect 262382 263218 262466 263454
rect 262702 263218 296146 263454
rect 296382 263218 296466 263454
rect 296702 263218 330146 263454
rect 330382 263218 330466 263454
rect 330702 263218 364146 263454
rect 364382 263218 364466 263454
rect 364702 263218 398146 263454
rect 398382 263218 398466 263454
rect 398702 263218 432146 263454
rect 432382 263218 432466 263454
rect 432702 263218 466146 263454
rect 466382 263218 466466 263454
rect 466702 263218 500146 263454
rect 500382 263218 500466 263454
rect 500702 263218 534146 263454
rect 534382 263218 534466 263454
rect 534702 263218 568146 263454
rect 568382 263218 568466 263454
rect 568702 263218 591102 263454
rect 591338 263218 591422 263454
rect 591658 263218 592650 263454
rect -8726 263186 592650 263218
rect -8726 260054 592650 260086
rect -8726 259818 -6774 260054
rect -6538 259818 -6454 260054
rect -6218 259818 20426 260054
rect 20662 259818 20746 260054
rect 20982 259818 54426 260054
rect 54662 259818 54746 260054
rect 54982 259818 88426 260054
rect 88662 259818 88746 260054
rect 88982 259818 122426 260054
rect 122662 259818 122746 260054
rect 122982 259818 156426 260054
rect 156662 259818 156746 260054
rect 156982 259818 190426 260054
rect 190662 259818 190746 260054
rect 190982 259818 224426 260054
rect 224662 259818 224746 260054
rect 224982 259818 258426 260054
rect 258662 259818 258746 260054
rect 258982 259818 292426 260054
rect 292662 259818 292746 260054
rect 292982 259818 326426 260054
rect 326662 259818 326746 260054
rect 326982 259818 360426 260054
rect 360662 259818 360746 260054
rect 360982 259818 394426 260054
rect 394662 259818 394746 260054
rect 394982 259818 428426 260054
rect 428662 259818 428746 260054
rect 428982 259818 462426 260054
rect 462662 259818 462746 260054
rect 462982 259818 496426 260054
rect 496662 259818 496746 260054
rect 496982 259818 530426 260054
rect 530662 259818 530746 260054
rect 530982 259818 564426 260054
rect 564662 259818 564746 260054
rect 564982 259818 590142 260054
rect 590378 259818 590462 260054
rect 590698 259818 592650 260054
rect -8726 259734 592650 259818
rect -8726 259498 -6774 259734
rect -6538 259498 -6454 259734
rect -6218 259498 20426 259734
rect 20662 259498 20746 259734
rect 20982 259498 54426 259734
rect 54662 259498 54746 259734
rect 54982 259498 88426 259734
rect 88662 259498 88746 259734
rect 88982 259498 122426 259734
rect 122662 259498 122746 259734
rect 122982 259498 156426 259734
rect 156662 259498 156746 259734
rect 156982 259498 190426 259734
rect 190662 259498 190746 259734
rect 190982 259498 224426 259734
rect 224662 259498 224746 259734
rect 224982 259498 258426 259734
rect 258662 259498 258746 259734
rect 258982 259498 292426 259734
rect 292662 259498 292746 259734
rect 292982 259498 326426 259734
rect 326662 259498 326746 259734
rect 326982 259498 360426 259734
rect 360662 259498 360746 259734
rect 360982 259498 394426 259734
rect 394662 259498 394746 259734
rect 394982 259498 428426 259734
rect 428662 259498 428746 259734
rect 428982 259498 462426 259734
rect 462662 259498 462746 259734
rect 462982 259498 496426 259734
rect 496662 259498 496746 259734
rect 496982 259498 530426 259734
rect 530662 259498 530746 259734
rect 530982 259498 564426 259734
rect 564662 259498 564746 259734
rect 564982 259498 590142 259734
rect 590378 259498 590462 259734
rect 590698 259498 592650 259734
rect -8726 259466 592650 259498
rect -8726 256334 592650 256366
rect -8726 256098 -5814 256334
rect -5578 256098 -5494 256334
rect -5258 256098 16706 256334
rect 16942 256098 17026 256334
rect 17262 256098 50706 256334
rect 50942 256098 51026 256334
rect 51262 256098 84706 256334
rect 84942 256098 85026 256334
rect 85262 256098 118706 256334
rect 118942 256098 119026 256334
rect 119262 256098 152706 256334
rect 152942 256098 153026 256334
rect 153262 256098 186706 256334
rect 186942 256098 187026 256334
rect 187262 256098 220706 256334
rect 220942 256098 221026 256334
rect 221262 256098 254706 256334
rect 254942 256098 255026 256334
rect 255262 256098 288706 256334
rect 288942 256098 289026 256334
rect 289262 256098 322706 256334
rect 322942 256098 323026 256334
rect 323262 256098 356706 256334
rect 356942 256098 357026 256334
rect 357262 256098 390706 256334
rect 390942 256098 391026 256334
rect 391262 256098 424706 256334
rect 424942 256098 425026 256334
rect 425262 256098 458706 256334
rect 458942 256098 459026 256334
rect 459262 256098 492706 256334
rect 492942 256098 493026 256334
rect 493262 256098 526706 256334
rect 526942 256098 527026 256334
rect 527262 256098 560706 256334
rect 560942 256098 561026 256334
rect 561262 256098 589182 256334
rect 589418 256098 589502 256334
rect 589738 256098 592650 256334
rect -8726 256014 592650 256098
rect -8726 255778 -5814 256014
rect -5578 255778 -5494 256014
rect -5258 255778 16706 256014
rect 16942 255778 17026 256014
rect 17262 255778 50706 256014
rect 50942 255778 51026 256014
rect 51262 255778 84706 256014
rect 84942 255778 85026 256014
rect 85262 255778 118706 256014
rect 118942 255778 119026 256014
rect 119262 255778 152706 256014
rect 152942 255778 153026 256014
rect 153262 255778 186706 256014
rect 186942 255778 187026 256014
rect 187262 255778 220706 256014
rect 220942 255778 221026 256014
rect 221262 255778 254706 256014
rect 254942 255778 255026 256014
rect 255262 255778 288706 256014
rect 288942 255778 289026 256014
rect 289262 255778 322706 256014
rect 322942 255778 323026 256014
rect 323262 255778 356706 256014
rect 356942 255778 357026 256014
rect 357262 255778 390706 256014
rect 390942 255778 391026 256014
rect 391262 255778 424706 256014
rect 424942 255778 425026 256014
rect 425262 255778 458706 256014
rect 458942 255778 459026 256014
rect 459262 255778 492706 256014
rect 492942 255778 493026 256014
rect 493262 255778 526706 256014
rect 526942 255778 527026 256014
rect 527262 255778 560706 256014
rect 560942 255778 561026 256014
rect 561262 255778 589182 256014
rect 589418 255778 589502 256014
rect 589738 255778 592650 256014
rect -8726 255746 592650 255778
rect -8726 252614 592650 252646
rect -8726 252378 -4854 252614
rect -4618 252378 -4534 252614
rect -4298 252378 12986 252614
rect 13222 252378 13306 252614
rect 13542 252378 46986 252614
rect 47222 252378 47306 252614
rect 47542 252378 80986 252614
rect 81222 252378 81306 252614
rect 81542 252378 114986 252614
rect 115222 252378 115306 252614
rect 115542 252378 148986 252614
rect 149222 252378 149306 252614
rect 149542 252378 182986 252614
rect 183222 252378 183306 252614
rect 183542 252378 216986 252614
rect 217222 252378 217306 252614
rect 217542 252378 250986 252614
rect 251222 252378 251306 252614
rect 251542 252378 284986 252614
rect 285222 252378 285306 252614
rect 285542 252378 318986 252614
rect 319222 252378 319306 252614
rect 319542 252378 352986 252614
rect 353222 252378 353306 252614
rect 353542 252378 386986 252614
rect 387222 252378 387306 252614
rect 387542 252378 420986 252614
rect 421222 252378 421306 252614
rect 421542 252378 454986 252614
rect 455222 252378 455306 252614
rect 455542 252378 488986 252614
rect 489222 252378 489306 252614
rect 489542 252378 522986 252614
rect 523222 252378 523306 252614
rect 523542 252378 556986 252614
rect 557222 252378 557306 252614
rect 557542 252378 588222 252614
rect 588458 252378 588542 252614
rect 588778 252378 592650 252614
rect -8726 252294 592650 252378
rect -8726 252058 -4854 252294
rect -4618 252058 -4534 252294
rect -4298 252058 12986 252294
rect 13222 252058 13306 252294
rect 13542 252058 46986 252294
rect 47222 252058 47306 252294
rect 47542 252058 80986 252294
rect 81222 252058 81306 252294
rect 81542 252058 114986 252294
rect 115222 252058 115306 252294
rect 115542 252058 148986 252294
rect 149222 252058 149306 252294
rect 149542 252058 182986 252294
rect 183222 252058 183306 252294
rect 183542 252058 216986 252294
rect 217222 252058 217306 252294
rect 217542 252058 250986 252294
rect 251222 252058 251306 252294
rect 251542 252058 284986 252294
rect 285222 252058 285306 252294
rect 285542 252058 318986 252294
rect 319222 252058 319306 252294
rect 319542 252058 352986 252294
rect 353222 252058 353306 252294
rect 353542 252058 386986 252294
rect 387222 252058 387306 252294
rect 387542 252058 420986 252294
rect 421222 252058 421306 252294
rect 421542 252058 454986 252294
rect 455222 252058 455306 252294
rect 455542 252058 488986 252294
rect 489222 252058 489306 252294
rect 489542 252058 522986 252294
rect 523222 252058 523306 252294
rect 523542 252058 556986 252294
rect 557222 252058 557306 252294
rect 557542 252058 588222 252294
rect 588458 252058 588542 252294
rect 588778 252058 592650 252294
rect -8726 252026 592650 252058
rect -8726 248894 592650 248926
rect -8726 248658 -3894 248894
rect -3658 248658 -3574 248894
rect -3338 248658 9266 248894
rect 9502 248658 9586 248894
rect 9822 248658 43266 248894
rect 43502 248658 43586 248894
rect 43822 248658 77266 248894
rect 77502 248658 77586 248894
rect 77822 248658 111266 248894
rect 111502 248658 111586 248894
rect 111822 248658 145266 248894
rect 145502 248658 145586 248894
rect 145822 248658 179266 248894
rect 179502 248658 179586 248894
rect 179822 248658 213266 248894
rect 213502 248658 213586 248894
rect 213822 248658 247266 248894
rect 247502 248658 247586 248894
rect 247822 248658 281266 248894
rect 281502 248658 281586 248894
rect 281822 248658 315266 248894
rect 315502 248658 315586 248894
rect 315822 248658 349266 248894
rect 349502 248658 349586 248894
rect 349822 248658 383266 248894
rect 383502 248658 383586 248894
rect 383822 248658 417266 248894
rect 417502 248658 417586 248894
rect 417822 248658 451266 248894
rect 451502 248658 451586 248894
rect 451822 248658 485266 248894
rect 485502 248658 485586 248894
rect 485822 248658 519266 248894
rect 519502 248658 519586 248894
rect 519822 248658 553266 248894
rect 553502 248658 553586 248894
rect 553822 248658 587262 248894
rect 587498 248658 587582 248894
rect 587818 248658 592650 248894
rect -8726 248574 592650 248658
rect -8726 248338 -3894 248574
rect -3658 248338 -3574 248574
rect -3338 248338 9266 248574
rect 9502 248338 9586 248574
rect 9822 248338 43266 248574
rect 43502 248338 43586 248574
rect 43822 248338 77266 248574
rect 77502 248338 77586 248574
rect 77822 248338 111266 248574
rect 111502 248338 111586 248574
rect 111822 248338 145266 248574
rect 145502 248338 145586 248574
rect 145822 248338 179266 248574
rect 179502 248338 179586 248574
rect 179822 248338 213266 248574
rect 213502 248338 213586 248574
rect 213822 248338 247266 248574
rect 247502 248338 247586 248574
rect 247822 248338 281266 248574
rect 281502 248338 281586 248574
rect 281822 248338 315266 248574
rect 315502 248338 315586 248574
rect 315822 248338 349266 248574
rect 349502 248338 349586 248574
rect 349822 248338 383266 248574
rect 383502 248338 383586 248574
rect 383822 248338 417266 248574
rect 417502 248338 417586 248574
rect 417822 248338 451266 248574
rect 451502 248338 451586 248574
rect 451822 248338 485266 248574
rect 485502 248338 485586 248574
rect 485822 248338 519266 248574
rect 519502 248338 519586 248574
rect 519822 248338 553266 248574
rect 553502 248338 553586 248574
rect 553822 248338 587262 248574
rect 587498 248338 587582 248574
rect 587818 248338 592650 248574
rect -8726 248306 592650 248338
rect -8726 245174 592650 245206
rect -8726 244938 -2934 245174
rect -2698 244938 -2614 245174
rect -2378 244938 5546 245174
rect 5782 244938 5866 245174
rect 6102 244938 39546 245174
rect 39782 244938 39866 245174
rect 40102 244938 73546 245174
rect 73782 244938 73866 245174
rect 74102 244938 107546 245174
rect 107782 244938 107866 245174
rect 108102 244938 141546 245174
rect 141782 244938 141866 245174
rect 142102 244938 175546 245174
rect 175782 244938 175866 245174
rect 176102 244938 209546 245174
rect 209782 244938 209866 245174
rect 210102 244938 243546 245174
rect 243782 244938 243866 245174
rect 244102 244938 277546 245174
rect 277782 244938 277866 245174
rect 278102 244938 311546 245174
rect 311782 244938 311866 245174
rect 312102 244938 345546 245174
rect 345782 244938 345866 245174
rect 346102 244938 379546 245174
rect 379782 244938 379866 245174
rect 380102 244938 413546 245174
rect 413782 244938 413866 245174
rect 414102 244938 447546 245174
rect 447782 244938 447866 245174
rect 448102 244938 481546 245174
rect 481782 244938 481866 245174
rect 482102 244938 515546 245174
rect 515782 244938 515866 245174
rect 516102 244938 549546 245174
rect 549782 244938 549866 245174
rect 550102 244938 586302 245174
rect 586538 244938 586622 245174
rect 586858 244938 592650 245174
rect -8726 244854 592650 244938
rect -8726 244618 -2934 244854
rect -2698 244618 -2614 244854
rect -2378 244618 5546 244854
rect 5782 244618 5866 244854
rect 6102 244618 39546 244854
rect 39782 244618 39866 244854
rect 40102 244618 73546 244854
rect 73782 244618 73866 244854
rect 74102 244618 107546 244854
rect 107782 244618 107866 244854
rect 108102 244618 141546 244854
rect 141782 244618 141866 244854
rect 142102 244618 175546 244854
rect 175782 244618 175866 244854
rect 176102 244618 209546 244854
rect 209782 244618 209866 244854
rect 210102 244618 243546 244854
rect 243782 244618 243866 244854
rect 244102 244618 277546 244854
rect 277782 244618 277866 244854
rect 278102 244618 311546 244854
rect 311782 244618 311866 244854
rect 312102 244618 345546 244854
rect 345782 244618 345866 244854
rect 346102 244618 379546 244854
rect 379782 244618 379866 244854
rect 380102 244618 413546 244854
rect 413782 244618 413866 244854
rect 414102 244618 447546 244854
rect 447782 244618 447866 244854
rect 448102 244618 481546 244854
rect 481782 244618 481866 244854
rect 482102 244618 515546 244854
rect 515782 244618 515866 244854
rect 516102 244618 549546 244854
rect 549782 244618 549866 244854
rect 550102 244618 586302 244854
rect 586538 244618 586622 244854
rect 586858 244618 592650 244854
rect -8726 244586 592650 244618
rect -8726 241454 592650 241486
rect -8726 241218 -1974 241454
rect -1738 241218 -1654 241454
rect -1418 241218 1826 241454
rect 2062 241218 2146 241454
rect 2382 241218 35826 241454
rect 36062 241218 36146 241454
rect 36382 241218 69826 241454
rect 70062 241218 70146 241454
rect 70382 241218 103826 241454
rect 104062 241218 104146 241454
rect 104382 241218 137826 241454
rect 138062 241218 138146 241454
rect 138382 241218 171826 241454
rect 172062 241218 172146 241454
rect 172382 241218 205826 241454
rect 206062 241218 206146 241454
rect 206382 241218 239826 241454
rect 240062 241218 240146 241454
rect 240382 241218 273826 241454
rect 274062 241218 274146 241454
rect 274382 241218 307826 241454
rect 308062 241218 308146 241454
rect 308382 241218 341826 241454
rect 342062 241218 342146 241454
rect 342382 241218 375826 241454
rect 376062 241218 376146 241454
rect 376382 241218 409826 241454
rect 410062 241218 410146 241454
rect 410382 241218 443826 241454
rect 444062 241218 444146 241454
rect 444382 241218 477826 241454
rect 478062 241218 478146 241454
rect 478382 241218 511826 241454
rect 512062 241218 512146 241454
rect 512382 241218 545826 241454
rect 546062 241218 546146 241454
rect 546382 241218 579826 241454
rect 580062 241218 580146 241454
rect 580382 241218 585342 241454
rect 585578 241218 585662 241454
rect 585898 241218 592650 241454
rect -8726 241134 592650 241218
rect -8726 240898 -1974 241134
rect -1738 240898 -1654 241134
rect -1418 240898 1826 241134
rect 2062 240898 2146 241134
rect 2382 240898 35826 241134
rect 36062 240898 36146 241134
rect 36382 240898 69826 241134
rect 70062 240898 70146 241134
rect 70382 240898 103826 241134
rect 104062 240898 104146 241134
rect 104382 240898 137826 241134
rect 138062 240898 138146 241134
rect 138382 240898 171826 241134
rect 172062 240898 172146 241134
rect 172382 240898 205826 241134
rect 206062 240898 206146 241134
rect 206382 240898 239826 241134
rect 240062 240898 240146 241134
rect 240382 240898 273826 241134
rect 274062 240898 274146 241134
rect 274382 240898 307826 241134
rect 308062 240898 308146 241134
rect 308382 240898 341826 241134
rect 342062 240898 342146 241134
rect 342382 240898 375826 241134
rect 376062 240898 376146 241134
rect 376382 240898 409826 241134
rect 410062 240898 410146 241134
rect 410382 240898 443826 241134
rect 444062 240898 444146 241134
rect 444382 240898 477826 241134
rect 478062 240898 478146 241134
rect 478382 240898 511826 241134
rect 512062 240898 512146 241134
rect 512382 240898 545826 241134
rect 546062 240898 546146 241134
rect 546382 240898 579826 241134
rect 580062 240898 580146 241134
rect 580382 240898 585342 241134
rect 585578 240898 585662 241134
rect 585898 240898 592650 241134
rect -8726 240866 592650 240898
rect -8726 233494 592650 233526
rect -8726 233258 -8694 233494
rect -8458 233258 -8374 233494
rect -8138 233258 27866 233494
rect 28102 233258 28186 233494
rect 28422 233258 61866 233494
rect 62102 233258 62186 233494
rect 62422 233258 95866 233494
rect 96102 233258 96186 233494
rect 96422 233258 129866 233494
rect 130102 233258 130186 233494
rect 130422 233258 163866 233494
rect 164102 233258 164186 233494
rect 164422 233258 197866 233494
rect 198102 233258 198186 233494
rect 198422 233258 231866 233494
rect 232102 233258 232186 233494
rect 232422 233258 265866 233494
rect 266102 233258 266186 233494
rect 266422 233258 299866 233494
rect 300102 233258 300186 233494
rect 300422 233258 333866 233494
rect 334102 233258 334186 233494
rect 334422 233258 367866 233494
rect 368102 233258 368186 233494
rect 368422 233258 401866 233494
rect 402102 233258 402186 233494
rect 402422 233258 435866 233494
rect 436102 233258 436186 233494
rect 436422 233258 469866 233494
rect 470102 233258 470186 233494
rect 470422 233258 503866 233494
rect 504102 233258 504186 233494
rect 504422 233258 537866 233494
rect 538102 233258 538186 233494
rect 538422 233258 571866 233494
rect 572102 233258 572186 233494
rect 572422 233258 592062 233494
rect 592298 233258 592382 233494
rect 592618 233258 592650 233494
rect -8726 233174 592650 233258
rect -8726 232938 -8694 233174
rect -8458 232938 -8374 233174
rect -8138 232938 27866 233174
rect 28102 232938 28186 233174
rect 28422 232938 61866 233174
rect 62102 232938 62186 233174
rect 62422 232938 95866 233174
rect 96102 232938 96186 233174
rect 96422 232938 129866 233174
rect 130102 232938 130186 233174
rect 130422 232938 163866 233174
rect 164102 232938 164186 233174
rect 164422 232938 197866 233174
rect 198102 232938 198186 233174
rect 198422 232938 231866 233174
rect 232102 232938 232186 233174
rect 232422 232938 265866 233174
rect 266102 232938 266186 233174
rect 266422 232938 299866 233174
rect 300102 232938 300186 233174
rect 300422 232938 333866 233174
rect 334102 232938 334186 233174
rect 334422 232938 367866 233174
rect 368102 232938 368186 233174
rect 368422 232938 401866 233174
rect 402102 232938 402186 233174
rect 402422 232938 435866 233174
rect 436102 232938 436186 233174
rect 436422 232938 469866 233174
rect 470102 232938 470186 233174
rect 470422 232938 503866 233174
rect 504102 232938 504186 233174
rect 504422 232938 537866 233174
rect 538102 232938 538186 233174
rect 538422 232938 571866 233174
rect 572102 232938 572186 233174
rect 572422 232938 592062 233174
rect 592298 232938 592382 233174
rect 592618 232938 592650 233174
rect -8726 232906 592650 232938
rect -8726 229774 592650 229806
rect -8726 229538 -7734 229774
rect -7498 229538 -7414 229774
rect -7178 229538 24146 229774
rect 24382 229538 24466 229774
rect 24702 229538 58146 229774
rect 58382 229538 58466 229774
rect 58702 229771 92146 229774
rect 58702 229538 65339 229771
rect -8726 229535 65339 229538
rect 65575 229535 65659 229771
rect 65895 229535 65979 229771
rect 66215 229535 66299 229771
rect 66535 229535 66619 229771
rect 66855 229535 66939 229771
rect 67175 229535 67259 229771
rect 67495 229535 67579 229771
rect 67815 229535 67899 229771
rect 68135 229535 68219 229771
rect 68455 229535 68539 229771
rect 68775 229535 68859 229771
rect 69095 229535 69179 229771
rect 69415 229535 69499 229771
rect 69735 229535 69819 229771
rect 70055 229538 92146 229771
rect 92382 229538 92466 229774
rect 92702 229538 126146 229774
rect 126382 229538 126466 229774
rect 126702 229538 160146 229774
rect 160382 229538 160466 229774
rect 160702 229538 194146 229774
rect 194382 229538 194466 229774
rect 194702 229538 228146 229774
rect 228382 229538 228466 229774
rect 228702 229538 262146 229774
rect 262382 229538 262466 229774
rect 262702 229538 296146 229774
rect 296382 229538 296466 229774
rect 296702 229538 330146 229774
rect 330382 229538 330466 229774
rect 330702 229538 364146 229774
rect 364382 229538 364466 229774
rect 364702 229538 398146 229774
rect 398382 229538 398466 229774
rect 398702 229538 432146 229774
rect 432382 229538 432466 229774
rect 432702 229538 466146 229774
rect 466382 229538 466466 229774
rect 466702 229538 500146 229774
rect 500382 229538 500466 229774
rect 500702 229538 534146 229774
rect 534382 229538 534466 229774
rect 534702 229538 568146 229774
rect 568382 229538 568466 229774
rect 568702 229538 591102 229774
rect 591338 229538 591422 229774
rect 591658 229538 592650 229774
rect 70055 229535 592650 229538
rect -8726 229454 592650 229535
rect -8726 229218 -7734 229454
rect -7498 229218 -7414 229454
rect -7178 229218 24146 229454
rect 24382 229218 24466 229454
rect 24702 229218 58146 229454
rect 58382 229218 58466 229454
rect 58702 229451 92146 229454
rect 58702 229218 65339 229451
rect -8726 229215 65339 229218
rect 65575 229215 65659 229451
rect 65895 229215 65979 229451
rect 66215 229215 66299 229451
rect 66535 229215 66619 229451
rect 66855 229215 66939 229451
rect 67175 229215 67259 229451
rect 67495 229215 67579 229451
rect 67815 229215 67899 229451
rect 68135 229215 68219 229451
rect 68455 229215 68539 229451
rect 68775 229215 68859 229451
rect 69095 229215 69179 229451
rect 69415 229215 69499 229451
rect 69735 229215 69819 229451
rect 70055 229218 92146 229451
rect 92382 229218 92466 229454
rect 92702 229218 126146 229454
rect 126382 229218 126466 229454
rect 126702 229218 160146 229454
rect 160382 229218 160466 229454
rect 160702 229218 194146 229454
rect 194382 229218 194466 229454
rect 194702 229218 228146 229454
rect 228382 229218 228466 229454
rect 228702 229218 262146 229454
rect 262382 229218 262466 229454
rect 262702 229218 296146 229454
rect 296382 229218 296466 229454
rect 296702 229218 330146 229454
rect 330382 229218 330466 229454
rect 330702 229218 364146 229454
rect 364382 229218 364466 229454
rect 364702 229218 398146 229454
rect 398382 229218 398466 229454
rect 398702 229218 432146 229454
rect 432382 229218 432466 229454
rect 432702 229218 466146 229454
rect 466382 229218 466466 229454
rect 466702 229218 500146 229454
rect 500382 229218 500466 229454
rect 500702 229218 534146 229454
rect 534382 229218 534466 229454
rect 534702 229218 568146 229454
rect 568382 229218 568466 229454
rect 568702 229218 591102 229454
rect 591338 229218 591422 229454
rect 591658 229218 592650 229454
rect 70055 229215 592650 229218
rect -8726 229186 592650 229215
rect -8726 226054 592650 226086
rect -8726 225818 -6774 226054
rect -6538 225818 -6454 226054
rect -6218 225818 20426 226054
rect 20662 225818 20746 226054
rect 20982 225991 190426 226054
rect 20982 225941 88426 225991
rect 20982 225818 54426 225941
rect -8726 225734 54426 225818
rect -8726 225498 -6774 225734
rect -6538 225498 -6454 225734
rect -6218 225498 20426 225734
rect 20662 225498 20746 225734
rect 20982 225705 54426 225734
rect 54662 225705 54746 225941
rect 54982 225801 88426 225941
rect 54982 225705 65462 225801
rect 20982 225565 65462 225705
rect 65698 225565 65782 225801
rect 66018 225565 66102 225801
rect 66338 225565 66422 225801
rect 66658 225565 66742 225801
rect 66978 225565 67062 225801
rect 67298 225565 67382 225801
rect 67618 225565 67702 225801
rect 67938 225565 68022 225801
rect 68258 225565 68342 225801
rect 68578 225565 68662 225801
rect 68898 225565 68982 225801
rect 69218 225565 69302 225801
rect 69538 225565 69622 225801
rect 69858 225565 69942 225801
rect 70178 225565 70262 225801
rect 70498 225565 70582 225801
rect 70818 225565 70902 225801
rect 71138 225755 88426 225801
rect 88662 225755 88746 225991
rect 88982 225755 122426 225991
rect 122662 225755 122746 225991
rect 122982 225755 156426 225991
rect 156662 225755 156746 225991
rect 156982 225818 190426 225991
rect 190662 225818 190746 226054
rect 190982 225991 428426 226054
rect 190982 225818 224426 225991
rect 156982 225755 224426 225818
rect 224662 225755 224746 225991
rect 224982 225755 258426 225991
rect 258662 225755 258746 225991
rect 258982 225755 292426 225991
rect 292662 225755 292746 225991
rect 292982 225755 326426 225991
rect 326662 225755 326746 225991
rect 326982 225755 360426 225991
rect 360662 225755 360746 225991
rect 360982 225755 394426 225991
rect 394662 225755 394746 225991
rect 394982 225818 428426 225991
rect 428662 225818 428746 226054
rect 428982 225818 462426 226054
rect 462662 225818 462746 226054
rect 462982 225818 496426 226054
rect 496662 225818 496746 226054
rect 496982 225818 530426 226054
rect 530662 225818 530746 226054
rect 530982 225818 564426 226054
rect 564662 225818 564746 226054
rect 564982 225818 590142 226054
rect 590378 225818 590462 226054
rect 590698 225818 592650 226054
rect 394982 225755 592650 225818
rect 71138 225734 592650 225755
rect 71138 225565 190426 225734
rect 20982 225498 190426 225565
rect 190662 225498 190746 225734
rect 190982 225498 428426 225734
rect 428662 225498 428746 225734
rect 428982 225498 462426 225734
rect 462662 225498 462746 225734
rect 462982 225498 496426 225734
rect 496662 225498 496746 225734
rect 496982 225498 530426 225734
rect 530662 225498 530746 225734
rect 530982 225498 564426 225734
rect 564662 225498 564746 225734
rect 564982 225498 590142 225734
rect 590378 225498 590462 225734
rect 590698 225498 592650 225734
rect -8726 225466 592650 225498
rect -8726 222334 592650 222366
rect -8726 222098 -5814 222334
rect -5578 222098 -5494 222334
rect -5258 222098 16706 222334
rect 16942 222098 17026 222334
rect 17262 222098 220706 222334
rect 220942 222098 221026 222334
rect 221262 222098 424706 222334
rect 424942 222098 425026 222334
rect 425262 222098 458706 222334
rect 458942 222098 459026 222334
rect 459262 222098 492706 222334
rect 492942 222098 493026 222334
rect 493262 222098 526706 222334
rect 526942 222098 527026 222334
rect 527262 222098 560706 222334
rect 560942 222098 561026 222334
rect 561262 222098 589182 222334
rect 589418 222098 589502 222334
rect 589738 222098 592650 222334
rect -8726 222014 592650 222098
rect -8726 221778 -5814 222014
rect -5578 221778 -5494 222014
rect -5258 221778 16706 222014
rect 16942 221778 17026 222014
rect 17262 221778 220706 222014
rect 220942 221778 221026 222014
rect 221262 221778 424706 222014
rect 424942 221778 425026 222014
rect 425262 221778 458706 222014
rect 458942 221778 459026 222014
rect 459262 221778 492706 222014
rect 492942 221778 493026 222014
rect 493262 221778 526706 222014
rect 526942 221778 527026 222014
rect 527262 221778 560706 222014
rect 560942 221778 561026 222014
rect 561262 221778 589182 222014
rect 589418 221778 589502 222014
rect 589738 221778 592650 222014
rect -8726 221746 592650 221778
rect -8726 218614 592650 218646
rect -8726 218378 -4854 218614
rect -4618 218378 -4534 218614
rect -4298 218378 12986 218614
rect 13222 218378 13306 218614
rect 13542 218378 250986 218614
rect 251222 218378 251306 218614
rect 251542 218378 420986 218614
rect 421222 218378 421306 218614
rect 421542 218378 454986 218614
rect 455222 218378 455306 218614
rect 455542 218378 488986 218614
rect 489222 218378 489306 218614
rect 489542 218378 522986 218614
rect 523222 218378 523306 218614
rect 523542 218378 556986 218614
rect 557222 218378 557306 218614
rect 557542 218378 588222 218614
rect 588458 218378 588542 218614
rect 588778 218378 592650 218614
rect -8726 218294 592650 218378
rect -8726 218058 -4854 218294
rect -4618 218058 -4534 218294
rect -4298 218058 12986 218294
rect 13222 218058 13306 218294
rect 13542 218058 250986 218294
rect 251222 218058 251306 218294
rect 251542 218058 420986 218294
rect 421222 218058 421306 218294
rect 421542 218058 454986 218294
rect 455222 218058 455306 218294
rect 455542 218058 488986 218294
rect 489222 218058 489306 218294
rect 489542 218058 522986 218294
rect 523222 218058 523306 218294
rect 523542 218058 556986 218294
rect 557222 218058 557306 218294
rect 557542 218058 588222 218294
rect 588458 218058 588542 218294
rect 588778 218058 592650 218294
rect -8726 218026 592650 218058
rect -8726 214894 592650 214926
rect -8726 214658 -3894 214894
rect -3658 214658 -3574 214894
rect -3338 214658 9266 214894
rect 9502 214658 9586 214894
rect 9822 214658 43266 214894
rect 43502 214658 43586 214894
rect 43822 214658 281266 214894
rect 281502 214658 281586 214894
rect 281822 214658 417266 214894
rect 417502 214658 417586 214894
rect 417822 214658 451266 214894
rect 451502 214658 451586 214894
rect 451822 214658 485266 214894
rect 485502 214658 485586 214894
rect 485822 214658 519266 214894
rect 519502 214658 519586 214894
rect 519822 214658 553266 214894
rect 553502 214658 553586 214894
rect 553822 214658 587262 214894
rect 587498 214658 587582 214894
rect 587818 214658 592650 214894
rect -8726 214574 592650 214658
rect -8726 214338 -3894 214574
rect -3658 214338 -3574 214574
rect -3338 214338 9266 214574
rect 9502 214338 9586 214574
rect 9822 214338 43266 214574
rect 43502 214338 43586 214574
rect 43822 214338 281266 214574
rect 281502 214338 281586 214574
rect 281822 214338 417266 214574
rect 417502 214338 417586 214574
rect 417822 214338 451266 214574
rect 451502 214338 451586 214574
rect 451822 214338 485266 214574
rect 485502 214338 485586 214574
rect 485822 214338 519266 214574
rect 519502 214338 519586 214574
rect 519822 214338 553266 214574
rect 553502 214338 553586 214574
rect 553822 214338 587262 214574
rect 587498 214338 587582 214574
rect 587818 214338 592650 214574
rect -8726 214306 592650 214338
rect -8726 211174 592650 211206
rect -8726 210938 -2934 211174
rect -2698 210938 -2614 211174
rect -2378 210938 5546 211174
rect 5782 210938 5866 211174
rect 6102 210938 39546 211174
rect 39782 210938 39866 211174
rect 40102 210938 73546 211174
rect 73782 210938 73866 211174
rect 74102 210938 107546 211174
rect 107782 210938 107866 211174
rect 108102 210938 175546 211174
rect 175782 210938 175866 211174
rect 176102 210938 209546 211174
rect 209782 210938 209866 211174
rect 210102 210938 243546 211174
rect 243782 210938 243866 211174
rect 244102 210938 277546 211174
rect 277782 210938 277866 211174
rect 278102 210938 311546 211174
rect 311782 210938 311866 211174
rect 312102 210938 345546 211174
rect 345782 210938 345866 211174
rect 346102 210938 379546 211174
rect 379782 210938 379866 211174
rect 380102 210938 413546 211174
rect 413782 210938 413866 211174
rect 414102 210938 447546 211174
rect 447782 210938 447866 211174
rect 448102 210938 481546 211174
rect 481782 210938 481866 211174
rect 482102 210938 515546 211174
rect 515782 210938 515866 211174
rect 516102 210938 549546 211174
rect 549782 210938 549866 211174
rect 550102 210938 586302 211174
rect 586538 210938 586622 211174
rect 586858 210938 592650 211174
rect -8726 210854 592650 210938
rect -8726 210618 -2934 210854
rect -2698 210618 -2614 210854
rect -2378 210618 5546 210854
rect 5782 210618 5866 210854
rect 6102 210618 39546 210854
rect 39782 210618 39866 210854
rect 40102 210618 73546 210854
rect 73782 210618 73866 210854
rect 74102 210618 107546 210854
rect 107782 210618 107866 210854
rect 108102 210618 175546 210854
rect 175782 210618 175866 210854
rect 176102 210618 209546 210854
rect 209782 210618 209866 210854
rect 210102 210618 243546 210854
rect 243782 210618 243866 210854
rect 244102 210618 277546 210854
rect 277782 210618 277866 210854
rect 278102 210618 311546 210854
rect 311782 210618 311866 210854
rect 312102 210618 345546 210854
rect 345782 210618 345866 210854
rect 346102 210618 379546 210854
rect 379782 210618 379866 210854
rect 380102 210618 413546 210854
rect 413782 210618 413866 210854
rect 414102 210618 447546 210854
rect 447782 210618 447866 210854
rect 448102 210618 481546 210854
rect 481782 210618 481866 210854
rect 482102 210618 515546 210854
rect 515782 210618 515866 210854
rect 516102 210618 549546 210854
rect 549782 210618 549866 210854
rect 550102 210618 586302 210854
rect 586538 210618 586622 210854
rect 586858 210618 592650 210854
rect -8726 210586 592650 210618
rect -8726 207454 592650 207486
rect -8726 207218 -1974 207454
rect -1738 207218 -1654 207454
rect -1418 207218 1826 207454
rect 2062 207218 2146 207454
rect 2382 207218 35826 207454
rect 36062 207218 36146 207454
rect 36382 207218 69826 207454
rect 70062 207218 70146 207454
rect 70382 207218 103826 207454
rect 104062 207218 104146 207454
rect 104382 207218 171826 207454
rect 172062 207218 172146 207454
rect 172382 207218 205826 207454
rect 206062 207218 206146 207454
rect 206382 207218 239826 207454
rect 240062 207218 240146 207454
rect 240382 207218 273826 207454
rect 274062 207218 274146 207454
rect 274382 207218 307826 207454
rect 308062 207218 308146 207454
rect 308382 207218 341826 207454
rect 342062 207218 342146 207454
rect 342382 207218 375826 207454
rect 376062 207218 376146 207454
rect 376382 207218 409826 207454
rect 410062 207218 410146 207454
rect 410382 207218 443826 207454
rect 444062 207218 444146 207454
rect 444382 207218 477826 207454
rect 478062 207218 478146 207454
rect 478382 207218 511826 207454
rect 512062 207218 512146 207454
rect 512382 207218 545826 207454
rect 546062 207218 546146 207454
rect 546382 207218 579826 207454
rect 580062 207218 580146 207454
rect 580382 207218 585342 207454
rect 585578 207218 585662 207454
rect 585898 207218 592650 207454
rect -8726 207134 592650 207218
rect -8726 206898 -1974 207134
rect -1738 206898 -1654 207134
rect -1418 206898 1826 207134
rect 2062 206898 2146 207134
rect 2382 206898 35826 207134
rect 36062 206898 36146 207134
rect 36382 206898 69826 207134
rect 70062 206898 70146 207134
rect 70382 206898 103826 207134
rect 104062 206898 104146 207134
rect 104382 206898 171826 207134
rect 172062 206898 172146 207134
rect 172382 206898 205826 207134
rect 206062 206898 206146 207134
rect 206382 206898 239826 207134
rect 240062 206898 240146 207134
rect 240382 206898 273826 207134
rect 274062 206898 274146 207134
rect 274382 206898 307826 207134
rect 308062 206898 308146 207134
rect 308382 206898 341826 207134
rect 342062 206898 342146 207134
rect 342382 206898 375826 207134
rect 376062 206898 376146 207134
rect 376382 206898 409826 207134
rect 410062 206898 410146 207134
rect 410382 206898 443826 207134
rect 444062 206898 444146 207134
rect 444382 206898 477826 207134
rect 478062 206898 478146 207134
rect 478382 206898 511826 207134
rect 512062 206898 512146 207134
rect 512382 206898 545826 207134
rect 546062 206898 546146 207134
rect 546382 206898 579826 207134
rect 580062 206898 580146 207134
rect 580382 206898 585342 207134
rect 585578 206898 585662 207134
rect 585898 206898 592650 207134
rect -8726 206866 592650 206898
rect -8726 199494 592650 199526
rect -8726 199258 -8694 199494
rect -8458 199258 -8374 199494
rect -8138 199258 27866 199494
rect 28102 199258 28186 199494
rect 28422 199258 61866 199494
rect 62102 199258 62186 199494
rect 62422 199258 95866 199494
rect 96102 199258 96186 199494
rect 96422 199258 129866 199494
rect 130102 199258 130186 199494
rect 130422 199258 163866 199494
rect 164102 199258 164186 199494
rect 164422 199258 197866 199494
rect 198102 199258 198186 199494
rect 198422 199258 231866 199494
rect 232102 199258 232186 199494
rect 232422 199258 265866 199494
rect 266102 199258 266186 199494
rect 266422 199258 299866 199494
rect 300102 199258 300186 199494
rect 300422 199258 333866 199494
rect 334102 199258 334186 199494
rect 334422 199258 367866 199494
rect 368102 199258 368186 199494
rect 368422 199258 401866 199494
rect 402102 199258 402186 199494
rect 402422 199258 435866 199494
rect 436102 199258 436186 199494
rect 436422 199258 469866 199494
rect 470102 199258 470186 199494
rect 470422 199258 503866 199494
rect 504102 199258 504186 199494
rect 504422 199258 537866 199494
rect 538102 199258 538186 199494
rect 538422 199258 571866 199494
rect 572102 199258 572186 199494
rect 572422 199258 592062 199494
rect 592298 199258 592382 199494
rect 592618 199258 592650 199494
rect -8726 199174 592650 199258
rect -8726 198938 -8694 199174
rect -8458 198938 -8374 199174
rect -8138 198938 27866 199174
rect 28102 198938 28186 199174
rect 28422 198938 61866 199174
rect 62102 198938 62186 199174
rect 62422 198938 95866 199174
rect 96102 198938 96186 199174
rect 96422 198938 129866 199174
rect 130102 198938 130186 199174
rect 130422 198938 163866 199174
rect 164102 198938 164186 199174
rect 164422 198938 197866 199174
rect 198102 198938 198186 199174
rect 198422 198938 231866 199174
rect 232102 198938 232186 199174
rect 232422 198938 265866 199174
rect 266102 198938 266186 199174
rect 266422 198938 299866 199174
rect 300102 198938 300186 199174
rect 300422 198938 333866 199174
rect 334102 198938 334186 199174
rect 334422 198938 367866 199174
rect 368102 198938 368186 199174
rect 368422 198938 401866 199174
rect 402102 198938 402186 199174
rect 402422 198938 435866 199174
rect 436102 198938 436186 199174
rect 436422 198938 469866 199174
rect 470102 198938 470186 199174
rect 470422 198938 503866 199174
rect 504102 198938 504186 199174
rect 504422 198938 537866 199174
rect 538102 198938 538186 199174
rect 538422 198938 571866 199174
rect 572102 198938 572186 199174
rect 572422 198938 592062 199174
rect 592298 198938 592382 199174
rect 592618 198938 592650 199174
rect -8726 198906 592650 198938
rect -8726 195774 592650 195806
rect -8726 195538 -7734 195774
rect -7498 195538 -7414 195774
rect -7178 195538 24146 195774
rect 24382 195538 24466 195774
rect 24702 195538 58146 195774
rect 58382 195538 58466 195774
rect 58702 195538 92146 195774
rect 92382 195538 92466 195774
rect 92702 195538 126146 195774
rect 126382 195538 126466 195774
rect 126702 195538 160146 195774
rect 160382 195538 160466 195774
rect 160702 195538 194146 195774
rect 194382 195538 194466 195774
rect 194702 195538 228146 195774
rect 228382 195538 228466 195774
rect 228702 195538 262146 195774
rect 262382 195538 262466 195774
rect 262702 195538 296146 195774
rect 296382 195538 296466 195774
rect 296702 195538 330146 195774
rect 330382 195538 330466 195774
rect 330702 195538 364146 195774
rect 364382 195538 364466 195774
rect 364702 195538 398146 195774
rect 398382 195538 398466 195774
rect 398702 195538 432146 195774
rect 432382 195538 432466 195774
rect 432702 195538 466146 195774
rect 466382 195538 466466 195774
rect 466702 195538 500146 195774
rect 500382 195538 500466 195774
rect 500702 195538 534146 195774
rect 534382 195538 534466 195774
rect 534702 195538 568146 195774
rect 568382 195538 568466 195774
rect 568702 195538 591102 195774
rect 591338 195538 591422 195774
rect 591658 195538 592650 195774
rect -8726 195454 592650 195538
rect -8726 195218 -7734 195454
rect -7498 195218 -7414 195454
rect -7178 195218 24146 195454
rect 24382 195218 24466 195454
rect 24702 195218 58146 195454
rect 58382 195218 58466 195454
rect 58702 195218 92146 195454
rect 92382 195218 92466 195454
rect 92702 195218 126146 195454
rect 126382 195218 126466 195454
rect 126702 195218 160146 195454
rect 160382 195218 160466 195454
rect 160702 195218 194146 195454
rect 194382 195218 194466 195454
rect 194702 195218 228146 195454
rect 228382 195218 228466 195454
rect 228702 195218 262146 195454
rect 262382 195218 262466 195454
rect 262702 195218 296146 195454
rect 296382 195218 296466 195454
rect 296702 195218 330146 195454
rect 330382 195218 330466 195454
rect 330702 195218 364146 195454
rect 364382 195218 364466 195454
rect 364702 195218 398146 195454
rect 398382 195218 398466 195454
rect 398702 195218 432146 195454
rect 432382 195218 432466 195454
rect 432702 195218 466146 195454
rect 466382 195218 466466 195454
rect 466702 195218 500146 195454
rect 500382 195218 500466 195454
rect 500702 195218 534146 195454
rect 534382 195218 534466 195454
rect 534702 195218 568146 195454
rect 568382 195218 568466 195454
rect 568702 195218 591102 195454
rect 591338 195218 591422 195454
rect 591658 195218 592650 195454
rect -8726 195186 592650 195218
rect -8726 192054 592650 192086
rect -8726 191818 -6774 192054
rect -6538 191818 -6454 192054
rect -6218 191818 20426 192054
rect 20662 191818 20746 192054
rect 20982 191818 54426 192054
rect 54662 191818 54746 192054
rect 54982 191818 88426 192054
rect 88662 191818 88746 192054
rect 88982 191818 122426 192054
rect 122662 191818 122746 192054
rect 122982 191818 190426 192054
rect 190662 191818 190746 192054
rect 190982 191818 224426 192054
rect 224662 191818 224746 192054
rect 224982 191818 258426 192054
rect 258662 191818 258746 192054
rect 258982 191818 292426 192054
rect 292662 191818 292746 192054
rect 292982 191818 326426 192054
rect 326662 191818 326746 192054
rect 326982 191818 360426 192054
rect 360662 191818 360746 192054
rect 360982 191818 394426 192054
rect 394662 191818 394746 192054
rect 394982 191818 428426 192054
rect 428662 191818 428746 192054
rect 428982 191818 462426 192054
rect 462662 191818 462746 192054
rect 462982 191818 496426 192054
rect 496662 191818 496746 192054
rect 496982 191818 530426 192054
rect 530662 191818 530746 192054
rect 530982 191818 564426 192054
rect 564662 191818 564746 192054
rect 564982 191818 590142 192054
rect 590378 191818 590462 192054
rect 590698 191818 592650 192054
rect -8726 191734 592650 191818
rect -8726 191498 -6774 191734
rect -6538 191498 -6454 191734
rect -6218 191498 20426 191734
rect 20662 191498 20746 191734
rect 20982 191498 54426 191734
rect 54662 191498 54746 191734
rect 54982 191498 88426 191734
rect 88662 191498 88746 191734
rect 88982 191498 122426 191734
rect 122662 191498 122746 191734
rect 122982 191498 190426 191734
rect 190662 191498 190746 191734
rect 190982 191498 224426 191734
rect 224662 191498 224746 191734
rect 224982 191498 258426 191734
rect 258662 191498 258746 191734
rect 258982 191498 292426 191734
rect 292662 191498 292746 191734
rect 292982 191498 326426 191734
rect 326662 191498 326746 191734
rect 326982 191498 360426 191734
rect 360662 191498 360746 191734
rect 360982 191498 394426 191734
rect 394662 191498 394746 191734
rect 394982 191498 428426 191734
rect 428662 191498 428746 191734
rect 428982 191498 462426 191734
rect 462662 191498 462746 191734
rect 462982 191498 496426 191734
rect 496662 191498 496746 191734
rect 496982 191498 530426 191734
rect 530662 191498 530746 191734
rect 530982 191498 564426 191734
rect 564662 191498 564746 191734
rect 564982 191498 590142 191734
rect 590378 191498 590462 191734
rect 590698 191498 592650 191734
rect -8726 191466 592650 191498
rect -8726 188334 592650 188366
rect -8726 188098 -5814 188334
rect -5578 188098 -5494 188334
rect -5258 188098 16706 188334
rect 16942 188098 17026 188334
rect 17262 188098 50706 188334
rect 50942 188098 51026 188334
rect 51262 188098 84706 188334
rect 84942 188098 85026 188334
rect 85262 188098 118706 188334
rect 118942 188098 119026 188334
rect 119262 188098 134376 188334
rect 134612 188098 134696 188334
rect 134932 188098 135016 188334
rect 135252 188098 135336 188334
rect 135572 188098 135656 188334
rect 135892 188098 135976 188334
rect 136212 188098 136296 188334
rect 136532 188098 136616 188334
rect 136852 188098 136936 188334
rect 137172 188098 137256 188334
rect 137492 188098 137576 188334
rect 137812 188098 137896 188334
rect 138132 188098 138216 188334
rect 138452 188098 138536 188334
rect 138772 188098 138856 188334
rect 139092 188098 139176 188334
rect 139412 188098 139496 188334
rect 139732 188098 139816 188334
rect 140052 188098 140136 188334
rect 140372 188098 140456 188334
rect 140692 188098 140776 188334
rect 141012 188098 141096 188334
rect 141332 188098 141416 188334
rect 141652 188098 141736 188334
rect 141972 188098 142056 188334
rect 142292 188098 142376 188334
rect 142612 188098 142696 188334
rect 142932 188098 143016 188334
rect 143252 188098 143336 188334
rect 143572 188098 143656 188334
rect 143892 188098 143976 188334
rect 144212 188098 144296 188334
rect 144532 188098 144616 188334
rect 144852 188098 144936 188334
rect 145172 188098 145256 188334
rect 145492 188098 145576 188334
rect 145812 188098 145896 188334
rect 146132 188098 146216 188334
rect 146452 188098 146536 188334
rect 146772 188098 146856 188334
rect 147092 188098 147176 188334
rect 147412 188098 147496 188334
rect 147732 188098 147816 188334
rect 148052 188098 148136 188334
rect 148372 188098 148456 188334
rect 148692 188098 148776 188334
rect 149012 188098 149096 188334
rect 149332 188098 149416 188334
rect 149652 188098 149736 188334
rect 149972 188098 150056 188334
rect 150292 188098 150376 188334
rect 150612 188098 150696 188334
rect 150932 188098 151016 188334
rect 151252 188098 151336 188334
rect 151572 188098 151656 188334
rect 151892 188098 151976 188334
rect 152212 188098 152296 188334
rect 152532 188098 152616 188334
rect 152852 188098 152936 188334
rect 153172 188098 153256 188334
rect 153492 188098 153576 188334
rect 153812 188098 153896 188334
rect 154132 188098 154216 188334
rect 154452 188098 154536 188334
rect 154772 188098 154856 188334
rect 155092 188098 155176 188334
rect 155412 188098 155496 188334
rect 155732 188098 155816 188334
rect 156052 188098 156136 188334
rect 156372 188098 156456 188334
rect 156692 188098 156776 188334
rect 157012 188098 157096 188334
rect 157332 188098 157416 188334
rect 157652 188098 157736 188334
rect 157972 188098 158056 188334
rect 158292 188098 158376 188334
rect 158612 188098 158696 188334
rect 158932 188098 159016 188334
rect 159252 188098 159336 188334
rect 159572 188098 159656 188334
rect 159892 188098 159976 188334
rect 160212 188098 160296 188334
rect 160532 188098 160616 188334
rect 160852 188098 160936 188334
rect 161172 188098 161256 188334
rect 161492 188098 161576 188334
rect 161812 188098 161896 188334
rect 162132 188098 162216 188334
rect 162452 188098 186706 188334
rect 186942 188098 187026 188334
rect 187262 188098 220706 188334
rect 220942 188098 221026 188334
rect 221262 188098 254706 188334
rect 254942 188098 255026 188334
rect 255262 188098 288706 188334
rect 288942 188098 289026 188334
rect 289262 188098 322706 188334
rect 322942 188098 323026 188334
rect 323262 188098 356706 188334
rect 356942 188098 357026 188334
rect 357262 188098 390706 188334
rect 390942 188098 391026 188334
rect 391262 188098 424706 188334
rect 424942 188098 425026 188334
rect 425262 188098 458706 188334
rect 458942 188098 459026 188334
rect 459262 188098 492706 188334
rect 492942 188098 493026 188334
rect 493262 188098 526706 188334
rect 526942 188098 527026 188334
rect 527262 188098 560706 188334
rect 560942 188098 561026 188334
rect 561262 188098 589182 188334
rect 589418 188098 589502 188334
rect 589738 188098 592650 188334
rect -8726 188014 592650 188098
rect -8726 187778 -5814 188014
rect -5578 187778 -5494 188014
rect -5258 187778 16706 188014
rect 16942 187778 17026 188014
rect 17262 187778 50706 188014
rect 50942 187778 51026 188014
rect 51262 187778 84706 188014
rect 84942 187778 85026 188014
rect 85262 187778 118706 188014
rect 118942 187778 119026 188014
rect 119262 187778 134376 188014
rect 134612 187778 134696 188014
rect 134932 187778 135016 188014
rect 135252 187778 135336 188014
rect 135572 187778 135656 188014
rect 135892 187778 135976 188014
rect 136212 187778 136296 188014
rect 136532 187778 136616 188014
rect 136852 187778 136936 188014
rect 137172 187778 137256 188014
rect 137492 187778 137576 188014
rect 137812 187778 137896 188014
rect 138132 187778 138216 188014
rect 138452 187778 138536 188014
rect 138772 187778 138856 188014
rect 139092 187778 139176 188014
rect 139412 187778 139496 188014
rect 139732 187778 139816 188014
rect 140052 187778 140136 188014
rect 140372 187778 140456 188014
rect 140692 187778 140776 188014
rect 141012 187778 141096 188014
rect 141332 187778 141416 188014
rect 141652 187778 141736 188014
rect 141972 187778 142056 188014
rect 142292 187778 142376 188014
rect 142612 187778 142696 188014
rect 142932 187778 143016 188014
rect 143252 187778 143336 188014
rect 143572 187778 143656 188014
rect 143892 187778 143976 188014
rect 144212 187778 144296 188014
rect 144532 187778 144616 188014
rect 144852 187778 144936 188014
rect 145172 187778 145256 188014
rect 145492 187778 145576 188014
rect 145812 187778 145896 188014
rect 146132 187778 146216 188014
rect 146452 187778 146536 188014
rect 146772 187778 146856 188014
rect 147092 187778 147176 188014
rect 147412 187778 147496 188014
rect 147732 187778 147816 188014
rect 148052 187778 148136 188014
rect 148372 187778 148456 188014
rect 148692 187778 148776 188014
rect 149012 187778 149096 188014
rect 149332 187778 149416 188014
rect 149652 187778 149736 188014
rect 149972 187778 150056 188014
rect 150292 187778 150376 188014
rect 150612 187778 150696 188014
rect 150932 187778 151016 188014
rect 151252 187778 151336 188014
rect 151572 187778 151656 188014
rect 151892 187778 151976 188014
rect 152212 187778 152296 188014
rect 152532 187778 152616 188014
rect 152852 187778 152936 188014
rect 153172 187778 153256 188014
rect 153492 187778 153576 188014
rect 153812 187778 153896 188014
rect 154132 187778 154216 188014
rect 154452 187778 154536 188014
rect 154772 187778 154856 188014
rect 155092 187778 155176 188014
rect 155412 187778 155496 188014
rect 155732 187778 155816 188014
rect 156052 187778 156136 188014
rect 156372 187778 156456 188014
rect 156692 187778 156776 188014
rect 157012 187778 157096 188014
rect 157332 187778 157416 188014
rect 157652 187778 157736 188014
rect 157972 187778 158056 188014
rect 158292 187778 158376 188014
rect 158612 187778 158696 188014
rect 158932 187778 159016 188014
rect 159252 187778 159336 188014
rect 159572 187778 159656 188014
rect 159892 187778 159976 188014
rect 160212 187778 160296 188014
rect 160532 187778 160616 188014
rect 160852 187778 160936 188014
rect 161172 187778 161256 188014
rect 161492 187778 161576 188014
rect 161812 187778 161896 188014
rect 162132 187778 162216 188014
rect 162452 187778 186706 188014
rect 186942 187778 187026 188014
rect 187262 187778 220706 188014
rect 220942 187778 221026 188014
rect 221262 187778 254706 188014
rect 254942 187778 255026 188014
rect 255262 187778 288706 188014
rect 288942 187778 289026 188014
rect 289262 187778 322706 188014
rect 322942 187778 323026 188014
rect 323262 187778 356706 188014
rect 356942 187778 357026 188014
rect 357262 187778 390706 188014
rect 390942 187778 391026 188014
rect 391262 187778 424706 188014
rect 424942 187778 425026 188014
rect 425262 187778 458706 188014
rect 458942 187778 459026 188014
rect 459262 187778 492706 188014
rect 492942 187778 493026 188014
rect 493262 187778 526706 188014
rect 526942 187778 527026 188014
rect 527262 187778 560706 188014
rect 560942 187778 561026 188014
rect 561262 187778 589182 188014
rect 589418 187778 589502 188014
rect 589738 187778 592650 188014
rect -8726 187746 592650 187778
rect -8726 184614 592650 184646
rect -8726 184378 -4854 184614
rect -4618 184378 -4534 184614
rect -4298 184378 12986 184614
rect 13222 184378 13306 184614
rect 13542 184378 46986 184614
rect 47222 184378 47306 184614
rect 47542 184378 80986 184614
rect 81222 184378 81306 184614
rect 81542 184378 114986 184614
rect 115222 184378 115306 184614
rect 115542 184378 148986 184614
rect 149222 184378 149306 184614
rect 149542 184378 182986 184614
rect 183222 184378 183306 184614
rect 183542 184378 216986 184614
rect 217222 184378 217306 184614
rect 217542 184378 250986 184614
rect 251222 184378 251306 184614
rect 251542 184378 284986 184614
rect 285222 184378 285306 184614
rect 285542 184378 318986 184614
rect 319222 184378 319306 184614
rect 319542 184378 352986 184614
rect 353222 184378 353306 184614
rect 353542 184378 386986 184614
rect 387222 184378 387306 184614
rect 387542 184378 420986 184614
rect 421222 184378 421306 184614
rect 421542 184378 454986 184614
rect 455222 184378 455306 184614
rect 455542 184378 488986 184614
rect 489222 184378 489306 184614
rect 489542 184378 522986 184614
rect 523222 184378 523306 184614
rect 523542 184378 556986 184614
rect 557222 184378 557306 184614
rect 557542 184378 588222 184614
rect 588458 184378 588542 184614
rect 588778 184378 592650 184614
rect -8726 184294 592650 184378
rect -8726 184058 -4854 184294
rect -4618 184058 -4534 184294
rect -4298 184058 12986 184294
rect 13222 184058 13306 184294
rect 13542 184058 46986 184294
rect 47222 184058 47306 184294
rect 47542 184058 80986 184294
rect 81222 184058 81306 184294
rect 81542 184058 114986 184294
rect 115222 184058 115306 184294
rect 115542 184058 148986 184294
rect 149222 184058 149306 184294
rect 149542 184058 182986 184294
rect 183222 184058 183306 184294
rect 183542 184058 216986 184294
rect 217222 184058 217306 184294
rect 217542 184058 250986 184294
rect 251222 184058 251306 184294
rect 251542 184058 284986 184294
rect 285222 184058 285306 184294
rect 285542 184058 318986 184294
rect 319222 184058 319306 184294
rect 319542 184058 352986 184294
rect 353222 184058 353306 184294
rect 353542 184058 386986 184294
rect 387222 184058 387306 184294
rect 387542 184058 420986 184294
rect 421222 184058 421306 184294
rect 421542 184058 454986 184294
rect 455222 184058 455306 184294
rect 455542 184058 488986 184294
rect 489222 184058 489306 184294
rect 489542 184058 522986 184294
rect 523222 184058 523306 184294
rect 523542 184058 556986 184294
rect 557222 184058 557306 184294
rect 557542 184058 588222 184294
rect 588458 184058 588542 184294
rect 588778 184058 592650 184294
rect -8726 184026 592650 184058
rect -8726 180894 592650 180926
rect -8726 180658 -3894 180894
rect -3658 180658 -3574 180894
rect -3338 180658 9266 180894
rect 9502 180658 9586 180894
rect 9822 180658 43266 180894
rect 43502 180658 43586 180894
rect 43822 180658 77266 180894
rect 77502 180658 77586 180894
rect 77822 180658 111266 180894
rect 111502 180658 111586 180894
rect 111822 180658 145266 180894
rect 145502 180658 145586 180894
rect 145822 180658 179266 180894
rect 179502 180658 179586 180894
rect 179822 180658 213266 180894
rect 213502 180658 213586 180894
rect 213822 180658 247266 180894
rect 247502 180658 247586 180894
rect 247822 180658 281266 180894
rect 281502 180658 281586 180894
rect 281822 180658 315266 180894
rect 315502 180658 315586 180894
rect 315822 180658 349266 180894
rect 349502 180658 349586 180894
rect 349822 180658 383266 180894
rect 383502 180658 383586 180894
rect 383822 180658 417266 180894
rect 417502 180658 417586 180894
rect 417822 180658 451266 180894
rect 451502 180658 451586 180894
rect 451822 180658 485266 180894
rect 485502 180658 485586 180894
rect 485822 180658 519266 180894
rect 519502 180658 519586 180894
rect 519822 180658 553266 180894
rect 553502 180658 553586 180894
rect 553822 180658 587262 180894
rect 587498 180658 587582 180894
rect 587818 180658 592650 180894
rect -8726 180574 592650 180658
rect -8726 180338 -3894 180574
rect -3658 180338 -3574 180574
rect -3338 180338 9266 180574
rect 9502 180338 9586 180574
rect 9822 180338 43266 180574
rect 43502 180338 43586 180574
rect 43822 180338 77266 180574
rect 77502 180338 77586 180574
rect 77822 180338 111266 180574
rect 111502 180338 111586 180574
rect 111822 180338 145266 180574
rect 145502 180338 145586 180574
rect 145822 180338 179266 180574
rect 179502 180338 179586 180574
rect 179822 180338 213266 180574
rect 213502 180338 213586 180574
rect 213822 180338 247266 180574
rect 247502 180338 247586 180574
rect 247822 180338 281266 180574
rect 281502 180338 281586 180574
rect 281822 180338 315266 180574
rect 315502 180338 315586 180574
rect 315822 180338 349266 180574
rect 349502 180338 349586 180574
rect 349822 180338 383266 180574
rect 383502 180338 383586 180574
rect 383822 180338 417266 180574
rect 417502 180338 417586 180574
rect 417822 180338 451266 180574
rect 451502 180338 451586 180574
rect 451822 180338 485266 180574
rect 485502 180338 485586 180574
rect 485822 180338 519266 180574
rect 519502 180338 519586 180574
rect 519822 180338 553266 180574
rect 553502 180338 553586 180574
rect 553822 180338 587262 180574
rect 587498 180338 587582 180574
rect 587818 180338 592650 180574
rect -8726 180306 592650 180338
rect -8726 177174 592650 177206
rect -8726 176938 -2934 177174
rect -2698 176938 -2614 177174
rect -2378 176938 5546 177174
rect 5782 176938 5866 177174
rect 6102 176938 39546 177174
rect 39782 176938 39866 177174
rect 40102 176938 73546 177174
rect 73782 176938 73866 177174
rect 74102 176938 107546 177174
rect 107782 176938 107866 177174
rect 108102 176938 175546 177174
rect 175782 176938 175866 177174
rect 176102 176938 209546 177174
rect 209782 176938 209866 177174
rect 210102 176938 243546 177174
rect 243782 176938 243866 177174
rect 244102 176938 277546 177174
rect 277782 176938 277866 177174
rect 278102 176938 311546 177174
rect 311782 176938 311866 177174
rect 312102 176938 345546 177174
rect 345782 176938 345866 177174
rect 346102 176938 379546 177174
rect 379782 176938 379866 177174
rect 380102 176938 413546 177174
rect 413782 176938 413866 177174
rect 414102 176938 447546 177174
rect 447782 176938 447866 177174
rect 448102 176938 481546 177174
rect 481782 176938 481866 177174
rect 482102 176938 515546 177174
rect 515782 176938 515866 177174
rect 516102 176938 549546 177174
rect 549782 176938 549866 177174
rect 550102 176938 586302 177174
rect 586538 176938 586622 177174
rect 586858 176938 592650 177174
rect -8726 176854 592650 176938
rect -8726 176618 -2934 176854
rect -2698 176618 -2614 176854
rect -2378 176618 5546 176854
rect 5782 176618 5866 176854
rect 6102 176618 39546 176854
rect 39782 176618 39866 176854
rect 40102 176618 73546 176854
rect 73782 176618 73866 176854
rect 74102 176618 107546 176854
rect 107782 176618 107866 176854
rect 108102 176618 175546 176854
rect 175782 176618 175866 176854
rect 176102 176618 209546 176854
rect 209782 176618 209866 176854
rect 210102 176618 243546 176854
rect 243782 176618 243866 176854
rect 244102 176618 277546 176854
rect 277782 176618 277866 176854
rect 278102 176618 311546 176854
rect 311782 176618 311866 176854
rect 312102 176618 345546 176854
rect 345782 176618 345866 176854
rect 346102 176618 379546 176854
rect 379782 176618 379866 176854
rect 380102 176618 413546 176854
rect 413782 176618 413866 176854
rect 414102 176618 447546 176854
rect 447782 176618 447866 176854
rect 448102 176618 481546 176854
rect 481782 176618 481866 176854
rect 482102 176618 515546 176854
rect 515782 176618 515866 176854
rect 516102 176618 549546 176854
rect 549782 176618 549866 176854
rect 550102 176618 586302 176854
rect 586538 176618 586622 176854
rect 586858 176618 592650 176854
rect -8726 176586 592650 176618
rect -8726 173454 592650 173486
rect -8726 173218 -1974 173454
rect -1738 173218 -1654 173454
rect -1418 173218 1826 173454
rect 2062 173218 2146 173454
rect 2382 173218 35826 173454
rect 36062 173218 36146 173454
rect 36382 173218 69826 173454
rect 70062 173218 70146 173454
rect 70382 173218 103826 173454
rect 104062 173218 104146 173454
rect 104382 173218 137826 173454
rect 138062 173218 138146 173454
rect 138382 173218 171826 173454
rect 172062 173218 172146 173454
rect 172382 173218 205826 173454
rect 206062 173218 206146 173454
rect 206382 173218 239826 173454
rect 240062 173218 240146 173454
rect 240382 173218 273826 173454
rect 274062 173218 274146 173454
rect 274382 173218 307826 173454
rect 308062 173218 308146 173454
rect 308382 173218 341826 173454
rect 342062 173218 342146 173454
rect 342382 173218 375826 173454
rect 376062 173218 376146 173454
rect 376382 173218 409826 173454
rect 410062 173218 410146 173454
rect 410382 173218 443826 173454
rect 444062 173218 444146 173454
rect 444382 173218 477826 173454
rect 478062 173218 478146 173454
rect 478382 173218 511826 173454
rect 512062 173218 512146 173454
rect 512382 173218 545826 173454
rect 546062 173218 546146 173454
rect 546382 173218 579826 173454
rect 580062 173218 580146 173454
rect 580382 173218 585342 173454
rect 585578 173218 585662 173454
rect 585898 173218 592650 173454
rect -8726 173134 592650 173218
rect -8726 172898 -1974 173134
rect -1738 172898 -1654 173134
rect -1418 172898 1826 173134
rect 2062 172898 2146 173134
rect 2382 172898 35826 173134
rect 36062 172898 36146 173134
rect 36382 172898 69826 173134
rect 70062 172898 70146 173134
rect 70382 172898 103826 173134
rect 104062 172898 104146 173134
rect 104382 172898 137826 173134
rect 138062 172898 138146 173134
rect 138382 172898 171826 173134
rect 172062 172898 172146 173134
rect 172382 172898 205826 173134
rect 206062 172898 206146 173134
rect 206382 172898 239826 173134
rect 240062 172898 240146 173134
rect 240382 172898 273826 173134
rect 274062 172898 274146 173134
rect 274382 172898 307826 173134
rect 308062 172898 308146 173134
rect 308382 172898 341826 173134
rect 342062 172898 342146 173134
rect 342382 172898 375826 173134
rect 376062 172898 376146 173134
rect 376382 172898 409826 173134
rect 410062 172898 410146 173134
rect 410382 172898 443826 173134
rect 444062 172898 444146 173134
rect 444382 172898 477826 173134
rect 478062 172898 478146 173134
rect 478382 172898 511826 173134
rect 512062 172898 512146 173134
rect 512382 172898 545826 173134
rect 546062 172898 546146 173134
rect 546382 172898 579826 173134
rect 580062 172898 580146 173134
rect 580382 172898 585342 173134
rect 585578 172898 585662 173134
rect 585898 172898 592650 173134
rect -8726 172866 592650 172898
rect -8726 165494 592650 165526
rect -8726 165258 -8694 165494
rect -8458 165258 -8374 165494
rect -8138 165258 27866 165494
rect 28102 165258 28186 165494
rect 28422 165258 61866 165494
rect 62102 165258 62186 165494
rect 62422 165258 95866 165494
rect 96102 165258 96186 165494
rect 96422 165258 129866 165494
rect 130102 165258 130186 165494
rect 130422 165258 163866 165494
rect 164102 165258 164186 165494
rect 164422 165258 197866 165494
rect 198102 165258 198186 165494
rect 198422 165258 231866 165494
rect 232102 165258 232186 165494
rect 232422 165258 265866 165494
rect 266102 165258 266186 165494
rect 266422 165258 299866 165494
rect 300102 165258 300186 165494
rect 300422 165258 333866 165494
rect 334102 165258 334186 165494
rect 334422 165258 367866 165494
rect 368102 165258 368186 165494
rect 368422 165258 401866 165494
rect 402102 165258 402186 165494
rect 402422 165258 435866 165494
rect 436102 165258 436186 165494
rect 436422 165258 469866 165494
rect 470102 165258 470186 165494
rect 470422 165258 503866 165494
rect 504102 165258 504186 165494
rect 504422 165258 537866 165494
rect 538102 165258 538186 165494
rect 538422 165258 571866 165494
rect 572102 165258 572186 165494
rect 572422 165258 592062 165494
rect 592298 165258 592382 165494
rect 592618 165258 592650 165494
rect -8726 165174 592650 165258
rect -8726 164938 -8694 165174
rect -8458 164938 -8374 165174
rect -8138 164938 27866 165174
rect 28102 164938 28186 165174
rect 28422 164938 61866 165174
rect 62102 164938 62186 165174
rect 62422 164938 95866 165174
rect 96102 164938 96186 165174
rect 96422 164938 129866 165174
rect 130102 164938 130186 165174
rect 130422 164938 163866 165174
rect 164102 164938 164186 165174
rect 164422 164938 197866 165174
rect 198102 164938 198186 165174
rect 198422 164938 231866 165174
rect 232102 164938 232186 165174
rect 232422 164938 265866 165174
rect 266102 164938 266186 165174
rect 266422 164938 299866 165174
rect 300102 164938 300186 165174
rect 300422 164938 333866 165174
rect 334102 164938 334186 165174
rect 334422 164938 367866 165174
rect 368102 164938 368186 165174
rect 368422 164938 401866 165174
rect 402102 164938 402186 165174
rect 402422 164938 435866 165174
rect 436102 164938 436186 165174
rect 436422 164938 469866 165174
rect 470102 164938 470186 165174
rect 470422 164938 503866 165174
rect 504102 164938 504186 165174
rect 504422 164938 537866 165174
rect 538102 164938 538186 165174
rect 538422 164938 571866 165174
rect 572102 164938 572186 165174
rect 572422 164938 592062 165174
rect 592298 164938 592382 165174
rect 592618 164938 592650 165174
rect -8726 164906 592650 164938
rect -8726 161781 592650 161806
rect -8726 161774 134446 161781
rect -8726 161538 -7734 161774
rect -7498 161538 -7414 161774
rect -7178 161538 24146 161774
rect 24382 161538 24466 161774
rect 24702 161538 58146 161774
rect 58382 161538 58466 161774
rect 58702 161538 92146 161774
rect 92382 161538 92466 161774
rect 92702 161538 126146 161774
rect 126382 161538 126466 161774
rect 126702 161545 134446 161774
rect 134682 161545 134766 161781
rect 135002 161774 592650 161781
rect 135002 161545 160146 161774
rect 126702 161538 160146 161545
rect 160382 161538 160466 161774
rect 160702 161538 194146 161774
rect 194382 161538 194466 161774
rect 194702 161538 228146 161774
rect 228382 161538 228466 161774
rect 228702 161538 262146 161774
rect 262382 161538 262466 161774
rect 262702 161538 296146 161774
rect 296382 161538 296466 161774
rect 296702 161538 330146 161774
rect 330382 161538 330466 161774
rect 330702 161538 364146 161774
rect 364382 161538 364466 161774
rect 364702 161538 398146 161774
rect 398382 161538 398466 161774
rect 398702 161538 432146 161774
rect 432382 161538 432466 161774
rect 432702 161538 466146 161774
rect 466382 161538 466466 161774
rect 466702 161538 500146 161774
rect 500382 161538 500466 161774
rect 500702 161538 534146 161774
rect 534382 161538 534466 161774
rect 534702 161538 568146 161774
rect 568382 161538 568466 161774
rect 568702 161538 591102 161774
rect 591338 161538 591422 161774
rect 591658 161538 592650 161774
rect -8726 161461 592650 161538
rect -8726 161454 134446 161461
rect -8726 161218 -7734 161454
rect -7498 161218 -7414 161454
rect -7178 161218 24146 161454
rect 24382 161218 24466 161454
rect 24702 161218 58146 161454
rect 58382 161218 58466 161454
rect 58702 161218 92146 161454
rect 92382 161218 92466 161454
rect 92702 161218 126146 161454
rect 126382 161218 126466 161454
rect 126702 161225 134446 161454
rect 134682 161225 134766 161461
rect 135002 161454 592650 161461
rect 135002 161225 160146 161454
rect 126702 161218 160146 161225
rect 160382 161218 160466 161454
rect 160702 161218 194146 161454
rect 194382 161218 194466 161454
rect 194702 161218 228146 161454
rect 228382 161218 228466 161454
rect 228702 161218 262146 161454
rect 262382 161218 262466 161454
rect 262702 161218 296146 161454
rect 296382 161218 296466 161454
rect 296702 161218 330146 161454
rect 330382 161218 330466 161454
rect 330702 161218 364146 161454
rect 364382 161218 364466 161454
rect 364702 161218 398146 161454
rect 398382 161218 398466 161454
rect 398702 161218 432146 161454
rect 432382 161218 432466 161454
rect 432702 161218 466146 161454
rect 466382 161218 466466 161454
rect 466702 161218 500146 161454
rect 500382 161218 500466 161454
rect 500702 161218 534146 161454
rect 534382 161218 534466 161454
rect 534702 161218 568146 161454
rect 568382 161218 568466 161454
rect 568702 161218 591102 161454
rect 591338 161218 591422 161454
rect 591658 161218 592650 161454
rect -8726 161186 592650 161218
rect -8726 158054 592650 158086
rect -8726 157818 -6774 158054
rect -6538 157818 -6454 158054
rect -6218 157818 20426 158054
rect 20662 157818 20746 158054
rect 20982 157818 54426 158054
rect 54662 157818 54746 158054
rect 54982 157818 88426 158054
rect 88662 157818 88746 158054
rect 88982 157818 122426 158054
rect 122662 157818 122746 158054
rect 122982 157818 190426 158054
rect 190662 157818 190746 158054
rect 190982 157818 224426 158054
rect 224662 157818 224746 158054
rect 224982 157818 258426 158054
rect 258662 157818 258746 158054
rect 258982 157818 292426 158054
rect 292662 157818 292746 158054
rect 292982 157818 326426 158054
rect 326662 157818 326746 158054
rect 326982 157818 360426 158054
rect 360662 157818 360746 158054
rect 360982 157818 394426 158054
rect 394662 157818 394746 158054
rect 394982 157818 428426 158054
rect 428662 157818 428746 158054
rect 428982 157818 462426 158054
rect 462662 157818 462746 158054
rect 462982 157818 496426 158054
rect 496662 157818 496746 158054
rect 496982 157818 530426 158054
rect 530662 157818 530746 158054
rect 530982 157818 564426 158054
rect 564662 157818 564746 158054
rect 564982 157818 590142 158054
rect 590378 157818 590462 158054
rect 590698 157818 592650 158054
rect -8726 157734 592650 157818
rect -8726 157498 -6774 157734
rect -6538 157498 -6454 157734
rect -6218 157498 20426 157734
rect 20662 157498 20746 157734
rect 20982 157498 54426 157734
rect 54662 157498 54746 157734
rect 54982 157498 88426 157734
rect 88662 157498 88746 157734
rect 88982 157498 122426 157734
rect 122662 157498 122746 157734
rect 122982 157498 190426 157734
rect 190662 157498 190746 157734
rect 190982 157498 224426 157734
rect 224662 157498 224746 157734
rect 224982 157498 258426 157734
rect 258662 157498 258746 157734
rect 258982 157498 292426 157734
rect 292662 157498 292746 157734
rect 292982 157498 326426 157734
rect 326662 157498 326746 157734
rect 326982 157498 360426 157734
rect 360662 157498 360746 157734
rect 360982 157498 394426 157734
rect 394662 157498 394746 157734
rect 394982 157498 428426 157734
rect 428662 157498 428746 157734
rect 428982 157498 462426 157734
rect 462662 157498 462746 157734
rect 462982 157498 496426 157734
rect 496662 157498 496746 157734
rect 496982 157498 530426 157734
rect 530662 157498 530746 157734
rect 530982 157498 564426 157734
rect 564662 157498 564746 157734
rect 564982 157498 590142 157734
rect 590378 157498 590462 157734
rect 590698 157498 592650 157734
rect -8726 157466 592650 157498
rect -8726 154334 592650 154366
rect -8726 154098 -5814 154334
rect -5578 154098 -5494 154334
rect -5258 154098 16706 154334
rect 16942 154098 17026 154334
rect 17262 154098 50706 154334
rect 50942 154098 51026 154334
rect 51262 154098 84706 154334
rect 84942 154098 85026 154334
rect 85262 154098 118706 154334
rect 118942 154098 119026 154334
rect 119262 154098 186706 154334
rect 186942 154098 187026 154334
rect 187262 154098 220706 154334
rect 220942 154098 221026 154334
rect 221262 154098 254706 154334
rect 254942 154098 255026 154334
rect 255262 154098 288706 154334
rect 288942 154098 289026 154334
rect 289262 154098 322706 154334
rect 322942 154098 323026 154334
rect 323262 154098 356706 154334
rect 356942 154098 357026 154334
rect 357262 154098 390706 154334
rect 390942 154098 391026 154334
rect 391262 154098 424706 154334
rect 424942 154098 425026 154334
rect 425262 154098 458706 154334
rect 458942 154098 459026 154334
rect 459262 154098 492706 154334
rect 492942 154098 493026 154334
rect 493262 154098 526706 154334
rect 526942 154098 527026 154334
rect 527262 154098 560706 154334
rect 560942 154098 561026 154334
rect 561262 154098 589182 154334
rect 589418 154098 589502 154334
rect 589738 154098 592650 154334
rect -8726 154014 592650 154098
rect -8726 153778 -5814 154014
rect -5578 153778 -5494 154014
rect -5258 153778 16706 154014
rect 16942 153778 17026 154014
rect 17262 153778 50706 154014
rect 50942 153778 51026 154014
rect 51262 153778 84706 154014
rect 84942 153778 85026 154014
rect 85262 153778 118706 154014
rect 118942 153778 119026 154014
rect 119262 153778 186706 154014
rect 186942 153778 187026 154014
rect 187262 153778 220706 154014
rect 220942 153778 221026 154014
rect 221262 153778 254706 154014
rect 254942 153778 255026 154014
rect 255262 153778 288706 154014
rect 288942 153778 289026 154014
rect 289262 153778 322706 154014
rect 322942 153778 323026 154014
rect 323262 153778 356706 154014
rect 356942 153778 357026 154014
rect 357262 153778 390706 154014
rect 390942 153778 391026 154014
rect 391262 153778 424706 154014
rect 424942 153778 425026 154014
rect 425262 153778 458706 154014
rect 458942 153778 459026 154014
rect 459262 153778 492706 154014
rect 492942 153778 493026 154014
rect 493262 153778 526706 154014
rect 526942 153778 527026 154014
rect 527262 153778 560706 154014
rect 560942 153778 561026 154014
rect 561262 153778 589182 154014
rect 589418 153778 589502 154014
rect 589738 153778 592650 154014
rect -8726 153746 592650 153778
rect -8726 150614 592650 150646
rect -8726 150378 -4854 150614
rect -4618 150378 -4534 150614
rect -4298 150378 12986 150614
rect 13222 150378 13306 150614
rect 13542 150378 46986 150614
rect 47222 150378 47306 150614
rect 47542 150378 80986 150614
rect 81222 150378 81306 150614
rect 81542 150378 114986 150614
rect 115222 150378 115306 150614
rect 115542 150378 182986 150614
rect 183222 150378 183306 150614
rect 183542 150378 216986 150614
rect 217222 150378 217306 150614
rect 217542 150378 250986 150614
rect 251222 150378 251306 150614
rect 251542 150378 284986 150614
rect 285222 150378 285306 150614
rect 285542 150378 318986 150614
rect 319222 150378 319306 150614
rect 319542 150378 352986 150614
rect 353222 150378 353306 150614
rect 353542 150378 386986 150614
rect 387222 150378 387306 150614
rect 387542 150378 420986 150614
rect 421222 150378 421306 150614
rect 421542 150378 454986 150614
rect 455222 150378 455306 150614
rect 455542 150378 488986 150614
rect 489222 150378 489306 150614
rect 489542 150378 522986 150614
rect 523222 150378 523306 150614
rect 523542 150378 556986 150614
rect 557222 150378 557306 150614
rect 557542 150378 588222 150614
rect 588458 150378 588542 150614
rect 588778 150378 592650 150614
rect -8726 150294 592650 150378
rect -8726 150058 -4854 150294
rect -4618 150058 -4534 150294
rect -4298 150058 12986 150294
rect 13222 150058 13306 150294
rect 13542 150058 46986 150294
rect 47222 150058 47306 150294
rect 47542 150058 80986 150294
rect 81222 150058 81306 150294
rect 81542 150058 114986 150294
rect 115222 150058 115306 150294
rect 115542 150058 182986 150294
rect 183222 150058 183306 150294
rect 183542 150058 216986 150294
rect 217222 150058 217306 150294
rect 217542 150058 250986 150294
rect 251222 150058 251306 150294
rect 251542 150058 284986 150294
rect 285222 150058 285306 150294
rect 285542 150058 318986 150294
rect 319222 150058 319306 150294
rect 319542 150058 352986 150294
rect 353222 150058 353306 150294
rect 353542 150058 386986 150294
rect 387222 150058 387306 150294
rect 387542 150058 420986 150294
rect 421222 150058 421306 150294
rect 421542 150058 454986 150294
rect 455222 150058 455306 150294
rect 455542 150058 488986 150294
rect 489222 150058 489306 150294
rect 489542 150058 522986 150294
rect 523222 150058 523306 150294
rect 523542 150058 556986 150294
rect 557222 150058 557306 150294
rect 557542 150058 588222 150294
rect 588458 150058 588542 150294
rect 588778 150058 592650 150294
rect -8726 150026 592650 150058
rect -8726 146894 592650 146926
rect -8726 146658 -3894 146894
rect -3658 146658 -3574 146894
rect -3338 146658 9266 146894
rect 9502 146658 9586 146894
rect 9822 146658 43266 146894
rect 43502 146658 43586 146894
rect 43822 146658 77266 146894
rect 77502 146658 77586 146894
rect 77822 146658 111266 146894
rect 111502 146658 111586 146894
rect 111822 146658 179266 146894
rect 179502 146658 179586 146894
rect 179822 146658 213266 146894
rect 213502 146658 213586 146894
rect 213822 146658 247266 146894
rect 247502 146658 247586 146894
rect 247822 146658 281266 146894
rect 281502 146658 281586 146894
rect 281822 146658 315266 146894
rect 315502 146658 315586 146894
rect 315822 146658 349266 146894
rect 349502 146658 349586 146894
rect 349822 146658 383266 146894
rect 383502 146658 383586 146894
rect 383822 146658 417266 146894
rect 417502 146658 417586 146894
rect 417822 146658 451266 146894
rect 451502 146658 451586 146894
rect 451822 146658 485266 146894
rect 485502 146658 485586 146894
rect 485822 146658 519266 146894
rect 519502 146658 519586 146894
rect 519822 146658 553266 146894
rect 553502 146658 553586 146894
rect 553822 146658 587262 146894
rect 587498 146658 587582 146894
rect 587818 146658 592650 146894
rect -8726 146574 592650 146658
rect -8726 146338 -3894 146574
rect -3658 146338 -3574 146574
rect -3338 146338 9266 146574
rect 9502 146338 9586 146574
rect 9822 146338 43266 146574
rect 43502 146338 43586 146574
rect 43822 146338 77266 146574
rect 77502 146338 77586 146574
rect 77822 146338 111266 146574
rect 111502 146338 111586 146574
rect 111822 146338 179266 146574
rect 179502 146338 179586 146574
rect 179822 146338 213266 146574
rect 213502 146338 213586 146574
rect 213822 146338 247266 146574
rect 247502 146338 247586 146574
rect 247822 146338 281266 146574
rect 281502 146338 281586 146574
rect 281822 146338 315266 146574
rect 315502 146338 315586 146574
rect 315822 146338 349266 146574
rect 349502 146338 349586 146574
rect 349822 146338 383266 146574
rect 383502 146338 383586 146574
rect 383822 146338 417266 146574
rect 417502 146338 417586 146574
rect 417822 146338 451266 146574
rect 451502 146338 451586 146574
rect 451822 146338 485266 146574
rect 485502 146338 485586 146574
rect 485822 146338 519266 146574
rect 519502 146338 519586 146574
rect 519822 146338 553266 146574
rect 553502 146338 553586 146574
rect 553822 146338 587262 146574
rect 587498 146338 587582 146574
rect 587818 146338 592650 146574
rect -8726 146306 592650 146338
rect -8726 143174 592650 143206
rect -8726 142938 -2934 143174
rect -2698 142938 -2614 143174
rect -2378 142938 5546 143174
rect 5782 142938 5866 143174
rect 6102 142938 39546 143174
rect 39782 142938 39866 143174
rect 40102 142938 73546 143174
rect 73782 142938 73866 143174
rect 74102 142938 107546 143174
rect 107782 142938 107866 143174
rect 108102 142938 175546 143174
rect 175782 142938 175866 143174
rect 176102 142938 209546 143174
rect 209782 142938 209866 143174
rect 210102 142938 243546 143174
rect 243782 142938 243866 143174
rect 244102 142938 277546 143174
rect 277782 142938 277866 143174
rect 278102 142938 311546 143174
rect 311782 142938 311866 143174
rect 312102 142938 345546 143174
rect 345782 142938 345866 143174
rect 346102 142938 379546 143174
rect 379782 142938 379866 143174
rect 380102 142938 413546 143174
rect 413782 142938 413866 143174
rect 414102 142938 447546 143174
rect 447782 142938 447866 143174
rect 448102 142938 481546 143174
rect 481782 142938 481866 143174
rect 482102 142938 515546 143174
rect 515782 142938 515866 143174
rect 516102 142938 549546 143174
rect 549782 142938 549866 143174
rect 550102 142938 586302 143174
rect 586538 142938 586622 143174
rect 586858 142938 592650 143174
rect -8726 142854 592650 142938
rect -8726 142618 -2934 142854
rect -2698 142618 -2614 142854
rect -2378 142618 5546 142854
rect 5782 142618 5866 142854
rect 6102 142618 39546 142854
rect 39782 142618 39866 142854
rect 40102 142618 73546 142854
rect 73782 142618 73866 142854
rect 74102 142618 107546 142854
rect 107782 142618 107866 142854
rect 108102 142618 175546 142854
rect 175782 142618 175866 142854
rect 176102 142618 209546 142854
rect 209782 142618 209866 142854
rect 210102 142618 243546 142854
rect 243782 142618 243866 142854
rect 244102 142618 277546 142854
rect 277782 142618 277866 142854
rect 278102 142618 311546 142854
rect 311782 142618 311866 142854
rect 312102 142618 345546 142854
rect 345782 142618 345866 142854
rect 346102 142618 379546 142854
rect 379782 142618 379866 142854
rect 380102 142618 413546 142854
rect 413782 142618 413866 142854
rect 414102 142618 447546 142854
rect 447782 142618 447866 142854
rect 448102 142618 481546 142854
rect 481782 142618 481866 142854
rect 482102 142618 515546 142854
rect 515782 142618 515866 142854
rect 516102 142618 549546 142854
rect 549782 142618 549866 142854
rect 550102 142618 586302 142854
rect 586538 142618 586622 142854
rect 586858 142618 592650 142854
rect -8726 142586 592650 142618
rect -8726 139454 592650 139486
rect -8726 139218 -1974 139454
rect -1738 139218 -1654 139454
rect -1418 139218 1826 139454
rect 2062 139218 2146 139454
rect 2382 139218 35826 139454
rect 36062 139218 36146 139454
rect 36382 139218 69826 139454
rect 70062 139218 70146 139454
rect 70382 139218 103826 139454
rect 104062 139218 104146 139454
rect 104382 139218 171826 139454
rect 172062 139218 172146 139454
rect 172382 139218 205826 139454
rect 206062 139218 206146 139454
rect 206382 139218 239826 139454
rect 240062 139218 240146 139454
rect 240382 139218 273826 139454
rect 274062 139218 274146 139454
rect 274382 139218 307826 139454
rect 308062 139218 308146 139454
rect 308382 139218 341826 139454
rect 342062 139218 342146 139454
rect 342382 139218 375826 139454
rect 376062 139218 376146 139454
rect 376382 139218 409826 139454
rect 410062 139218 410146 139454
rect 410382 139218 443826 139454
rect 444062 139218 444146 139454
rect 444382 139218 477826 139454
rect 478062 139218 478146 139454
rect 478382 139218 511826 139454
rect 512062 139218 512146 139454
rect 512382 139218 545826 139454
rect 546062 139218 546146 139454
rect 546382 139218 579826 139454
rect 580062 139218 580146 139454
rect 580382 139218 585342 139454
rect 585578 139218 585662 139454
rect 585898 139218 592650 139454
rect -8726 139134 592650 139218
rect -8726 138898 -1974 139134
rect -1738 138898 -1654 139134
rect -1418 138898 1826 139134
rect 2062 138898 2146 139134
rect 2382 138898 35826 139134
rect 36062 138898 36146 139134
rect 36382 138898 69826 139134
rect 70062 138898 70146 139134
rect 70382 138898 103826 139134
rect 104062 138898 104146 139134
rect 104382 138898 171826 139134
rect 172062 138898 172146 139134
rect 172382 138898 205826 139134
rect 206062 138898 206146 139134
rect 206382 138898 239826 139134
rect 240062 138898 240146 139134
rect 240382 138898 273826 139134
rect 274062 138898 274146 139134
rect 274382 138898 307826 139134
rect 308062 138898 308146 139134
rect 308382 138898 341826 139134
rect 342062 138898 342146 139134
rect 342382 138898 375826 139134
rect 376062 138898 376146 139134
rect 376382 138898 409826 139134
rect 410062 138898 410146 139134
rect 410382 138898 443826 139134
rect 444062 138898 444146 139134
rect 444382 138898 477826 139134
rect 478062 138898 478146 139134
rect 478382 138898 511826 139134
rect 512062 138898 512146 139134
rect 512382 138898 545826 139134
rect 546062 138898 546146 139134
rect 546382 138898 579826 139134
rect 580062 138898 580146 139134
rect 580382 138898 585342 139134
rect 585578 138898 585662 139134
rect 585898 138898 592650 139134
rect -8726 138866 592650 138898
rect -8726 131494 592650 131526
rect -8726 131258 -8694 131494
rect -8458 131258 -8374 131494
rect -8138 131258 27866 131494
rect 28102 131258 28186 131494
rect 28422 131258 61866 131494
rect 62102 131258 62186 131494
rect 62422 131258 95866 131494
rect 96102 131258 96186 131494
rect 96422 131258 197866 131494
rect 198102 131258 198186 131494
rect 198422 131258 231866 131494
rect 232102 131258 232186 131494
rect 232422 131258 265866 131494
rect 266102 131258 266186 131494
rect 266422 131258 299866 131494
rect 300102 131258 300186 131494
rect 300422 131258 333866 131494
rect 334102 131258 334186 131494
rect 334422 131258 367866 131494
rect 368102 131258 368186 131494
rect 368422 131258 401866 131494
rect 402102 131258 402186 131494
rect 402422 131258 435866 131494
rect 436102 131258 436186 131494
rect 436422 131258 469866 131494
rect 470102 131258 470186 131494
rect 470422 131258 503866 131494
rect 504102 131258 504186 131494
rect 504422 131258 537866 131494
rect 538102 131258 538186 131494
rect 538422 131258 571866 131494
rect 572102 131258 572186 131494
rect 572422 131258 592062 131494
rect 592298 131258 592382 131494
rect 592618 131258 592650 131494
rect -8726 131174 592650 131258
rect -8726 130938 -8694 131174
rect -8458 130938 -8374 131174
rect -8138 130938 27866 131174
rect 28102 130938 28186 131174
rect 28422 130938 61866 131174
rect 62102 130938 62186 131174
rect 62422 130938 95866 131174
rect 96102 130938 96186 131174
rect 96422 130938 197866 131174
rect 198102 130938 198186 131174
rect 198422 130938 231866 131174
rect 232102 130938 232186 131174
rect 232422 130938 265866 131174
rect 266102 130938 266186 131174
rect 266422 130938 299866 131174
rect 300102 130938 300186 131174
rect 300422 130938 333866 131174
rect 334102 130938 334186 131174
rect 334422 130938 367866 131174
rect 368102 130938 368186 131174
rect 368422 130938 401866 131174
rect 402102 130938 402186 131174
rect 402422 130938 435866 131174
rect 436102 130938 436186 131174
rect 436422 130938 469866 131174
rect 470102 130938 470186 131174
rect 470422 130938 503866 131174
rect 504102 130938 504186 131174
rect 504422 130938 537866 131174
rect 538102 130938 538186 131174
rect 538422 130938 571866 131174
rect 572102 130938 572186 131174
rect 572422 130938 592062 131174
rect 592298 130938 592382 131174
rect 592618 130938 592650 131174
rect -8726 130906 592650 130938
rect -8726 127774 592650 127806
rect -8726 127538 -7734 127774
rect -7498 127538 -7414 127774
rect -7178 127538 24146 127774
rect 24382 127538 24466 127774
rect 24702 127538 58146 127774
rect 58382 127538 58466 127774
rect 58702 127538 92146 127774
rect 92382 127538 92466 127774
rect 92702 127538 194146 127774
rect 194382 127538 194466 127774
rect 194702 127538 228146 127774
rect 228382 127538 228466 127774
rect 228702 127538 262146 127774
rect 262382 127538 262466 127774
rect 262702 127538 296146 127774
rect 296382 127538 296466 127774
rect 296702 127538 330146 127774
rect 330382 127538 330466 127774
rect 330702 127538 364146 127774
rect 364382 127538 364466 127774
rect 364702 127538 398146 127774
rect 398382 127538 398466 127774
rect 398702 127538 432146 127774
rect 432382 127538 432466 127774
rect 432702 127538 466146 127774
rect 466382 127538 466466 127774
rect 466702 127538 500146 127774
rect 500382 127538 500466 127774
rect 500702 127538 534146 127774
rect 534382 127538 534466 127774
rect 534702 127538 568146 127774
rect 568382 127538 568466 127774
rect 568702 127538 591102 127774
rect 591338 127538 591422 127774
rect 591658 127538 592650 127774
rect -8726 127454 592650 127538
rect -8726 127218 -7734 127454
rect -7498 127218 -7414 127454
rect -7178 127218 24146 127454
rect 24382 127218 24466 127454
rect 24702 127218 58146 127454
rect 58382 127218 58466 127454
rect 58702 127218 92146 127454
rect 92382 127218 92466 127454
rect 92702 127218 194146 127454
rect 194382 127218 194466 127454
rect 194702 127218 228146 127454
rect 228382 127218 228466 127454
rect 228702 127218 262146 127454
rect 262382 127218 262466 127454
rect 262702 127218 296146 127454
rect 296382 127218 296466 127454
rect 296702 127218 330146 127454
rect 330382 127218 330466 127454
rect 330702 127218 364146 127454
rect 364382 127218 364466 127454
rect 364702 127218 398146 127454
rect 398382 127218 398466 127454
rect 398702 127218 432146 127454
rect 432382 127218 432466 127454
rect 432702 127218 466146 127454
rect 466382 127218 466466 127454
rect 466702 127218 500146 127454
rect 500382 127218 500466 127454
rect 500702 127218 534146 127454
rect 534382 127218 534466 127454
rect 534702 127218 568146 127454
rect 568382 127218 568466 127454
rect 568702 127218 591102 127454
rect 591338 127218 591422 127454
rect 591658 127218 592650 127454
rect -8726 127186 592650 127218
rect -8726 124054 592650 124086
rect -8726 123818 -6774 124054
rect -6538 123818 -6454 124054
rect -6218 123818 20426 124054
rect 20662 123818 20746 124054
rect 20982 123818 54426 124054
rect 54662 123818 54746 124054
rect 54982 123818 88426 124054
rect 88662 123818 88746 124054
rect 88982 123818 190426 124054
rect 190662 123818 190746 124054
rect 190982 123818 224426 124054
rect 224662 123818 224746 124054
rect 224982 123818 258426 124054
rect 258662 123818 258746 124054
rect 258982 123818 292426 124054
rect 292662 123818 292746 124054
rect 292982 123818 326426 124054
rect 326662 123818 326746 124054
rect 326982 123818 360426 124054
rect 360662 123818 360746 124054
rect 360982 123818 394426 124054
rect 394662 123818 394746 124054
rect 394982 123818 428426 124054
rect 428662 123818 428746 124054
rect 428982 123818 462426 124054
rect 462662 123818 462746 124054
rect 462982 123818 496426 124054
rect 496662 123818 496746 124054
rect 496982 123818 530426 124054
rect 530662 123818 530746 124054
rect 530982 123818 564426 124054
rect 564662 123818 564746 124054
rect 564982 123818 590142 124054
rect 590378 123818 590462 124054
rect 590698 123818 592650 124054
rect -8726 123734 592650 123818
rect -8726 123498 -6774 123734
rect -6538 123498 -6454 123734
rect -6218 123498 20426 123734
rect 20662 123498 20746 123734
rect 20982 123498 54426 123734
rect 54662 123498 54746 123734
rect 54982 123498 88426 123734
rect 88662 123498 88746 123734
rect 88982 123498 190426 123734
rect 190662 123498 190746 123734
rect 190982 123498 224426 123734
rect 224662 123498 224746 123734
rect 224982 123498 258426 123734
rect 258662 123498 258746 123734
rect 258982 123498 292426 123734
rect 292662 123498 292746 123734
rect 292982 123498 326426 123734
rect 326662 123498 326746 123734
rect 326982 123498 360426 123734
rect 360662 123498 360746 123734
rect 360982 123498 394426 123734
rect 394662 123498 394746 123734
rect 394982 123498 428426 123734
rect 428662 123498 428746 123734
rect 428982 123498 462426 123734
rect 462662 123498 462746 123734
rect 462982 123498 496426 123734
rect 496662 123498 496746 123734
rect 496982 123498 530426 123734
rect 530662 123498 530746 123734
rect 530982 123498 564426 123734
rect 564662 123498 564746 123734
rect 564982 123498 590142 123734
rect 590378 123498 590462 123734
rect 590698 123498 592650 123734
rect -8726 123466 592650 123498
rect -8726 120334 592650 120366
rect -8726 120098 -5814 120334
rect -5578 120098 -5494 120334
rect -5258 120098 16706 120334
rect 16942 120098 17026 120334
rect 17262 120098 50706 120334
rect 50942 120098 51026 120334
rect 51262 120098 84706 120334
rect 84942 120098 85026 120334
rect 85262 120098 186706 120334
rect 186942 120098 187026 120334
rect 187262 120098 220706 120334
rect 220942 120098 221026 120334
rect 221262 120098 254706 120334
rect 254942 120098 255026 120334
rect 255262 120098 288706 120334
rect 288942 120098 289026 120334
rect 289262 120098 322706 120334
rect 322942 120098 323026 120334
rect 323262 120098 356706 120334
rect 356942 120098 357026 120334
rect 357262 120098 390706 120334
rect 390942 120098 391026 120334
rect 391262 120098 424706 120334
rect 424942 120098 425026 120334
rect 425262 120098 458706 120334
rect 458942 120098 459026 120334
rect 459262 120098 492706 120334
rect 492942 120098 493026 120334
rect 493262 120098 526706 120334
rect 526942 120098 527026 120334
rect 527262 120098 560706 120334
rect 560942 120098 561026 120334
rect 561262 120098 589182 120334
rect 589418 120098 589502 120334
rect 589738 120098 592650 120334
rect -8726 120014 592650 120098
rect -8726 119778 -5814 120014
rect -5578 119778 -5494 120014
rect -5258 119778 16706 120014
rect 16942 119778 17026 120014
rect 17262 119778 50706 120014
rect 50942 119778 51026 120014
rect 51262 119778 84706 120014
rect 84942 119778 85026 120014
rect 85262 119778 186706 120014
rect 186942 119778 187026 120014
rect 187262 119778 220706 120014
rect 220942 119778 221026 120014
rect 221262 119778 254706 120014
rect 254942 119778 255026 120014
rect 255262 119778 288706 120014
rect 288942 119778 289026 120014
rect 289262 119778 322706 120014
rect 322942 119778 323026 120014
rect 323262 119778 356706 120014
rect 356942 119778 357026 120014
rect 357262 119778 390706 120014
rect 390942 119778 391026 120014
rect 391262 119778 424706 120014
rect 424942 119778 425026 120014
rect 425262 119778 458706 120014
rect 458942 119778 459026 120014
rect 459262 119778 492706 120014
rect 492942 119778 493026 120014
rect 493262 119778 526706 120014
rect 526942 119778 527026 120014
rect 527262 119778 560706 120014
rect 560942 119778 561026 120014
rect 561262 119778 589182 120014
rect 589418 119778 589502 120014
rect 589738 119778 592650 120014
rect -8726 119746 592650 119778
rect -8726 116614 592650 116646
rect -8726 116378 -4854 116614
rect -4618 116378 -4534 116614
rect -4298 116378 12986 116614
rect 13222 116378 13306 116614
rect 13542 116378 46986 116614
rect 47222 116378 47306 116614
rect 47542 116378 80986 116614
rect 81222 116378 81306 116614
rect 81542 116378 114986 116614
rect 115222 116378 115306 116614
rect 115542 116378 182986 116614
rect 183222 116378 183306 116614
rect 183542 116378 216986 116614
rect 217222 116378 217306 116614
rect 217542 116378 250986 116614
rect 251222 116378 251306 116614
rect 251542 116378 284986 116614
rect 285222 116378 285306 116614
rect 285542 116378 318986 116614
rect 319222 116378 319306 116614
rect 319542 116378 352986 116614
rect 353222 116378 353306 116614
rect 353542 116378 386986 116614
rect 387222 116378 387306 116614
rect 387542 116378 420986 116614
rect 421222 116378 421306 116614
rect 421542 116378 454986 116614
rect 455222 116378 455306 116614
rect 455542 116378 488986 116614
rect 489222 116378 489306 116614
rect 489542 116378 522986 116614
rect 523222 116378 523306 116614
rect 523542 116378 556986 116614
rect 557222 116378 557306 116614
rect 557542 116378 588222 116614
rect 588458 116378 588542 116614
rect 588778 116378 592650 116614
rect -8726 116294 592650 116378
rect -8726 116058 -4854 116294
rect -4618 116058 -4534 116294
rect -4298 116058 12986 116294
rect 13222 116058 13306 116294
rect 13542 116058 46986 116294
rect 47222 116058 47306 116294
rect 47542 116058 80986 116294
rect 81222 116058 81306 116294
rect 81542 116058 114986 116294
rect 115222 116058 115306 116294
rect 115542 116058 182986 116294
rect 183222 116058 183306 116294
rect 183542 116058 216986 116294
rect 217222 116058 217306 116294
rect 217542 116058 250986 116294
rect 251222 116058 251306 116294
rect 251542 116058 284986 116294
rect 285222 116058 285306 116294
rect 285542 116058 318986 116294
rect 319222 116058 319306 116294
rect 319542 116058 352986 116294
rect 353222 116058 353306 116294
rect 353542 116058 386986 116294
rect 387222 116058 387306 116294
rect 387542 116058 420986 116294
rect 421222 116058 421306 116294
rect 421542 116058 454986 116294
rect 455222 116058 455306 116294
rect 455542 116058 488986 116294
rect 489222 116058 489306 116294
rect 489542 116058 522986 116294
rect 523222 116058 523306 116294
rect 523542 116058 556986 116294
rect 557222 116058 557306 116294
rect 557542 116058 588222 116294
rect 588458 116058 588542 116294
rect 588778 116058 592650 116294
rect -8726 116026 592650 116058
rect -8726 112894 592650 112926
rect -8726 112658 -3894 112894
rect -3658 112658 -3574 112894
rect -3338 112658 9266 112894
rect 9502 112658 9586 112894
rect 9822 112658 43266 112894
rect 43502 112658 43586 112894
rect 43822 112658 77266 112894
rect 77502 112658 77586 112894
rect 77822 112658 111266 112894
rect 111502 112658 111586 112894
rect 111822 112658 179266 112894
rect 179502 112658 179586 112894
rect 179822 112658 213266 112894
rect 213502 112658 213586 112894
rect 213822 112658 247266 112894
rect 247502 112658 247586 112894
rect 247822 112658 281266 112894
rect 281502 112658 281586 112894
rect 281822 112658 315266 112894
rect 315502 112658 315586 112894
rect 315822 112658 349266 112894
rect 349502 112658 349586 112894
rect 349822 112658 383266 112894
rect 383502 112658 383586 112894
rect 383822 112658 417266 112894
rect 417502 112658 417586 112894
rect 417822 112658 451266 112894
rect 451502 112658 451586 112894
rect 451822 112658 485266 112894
rect 485502 112658 485586 112894
rect 485822 112658 519266 112894
rect 519502 112658 519586 112894
rect 519822 112658 553266 112894
rect 553502 112658 553586 112894
rect 553822 112658 587262 112894
rect 587498 112658 587582 112894
rect 587818 112658 592650 112894
rect -8726 112574 592650 112658
rect -8726 112338 -3894 112574
rect -3658 112338 -3574 112574
rect -3338 112338 9266 112574
rect 9502 112338 9586 112574
rect 9822 112338 43266 112574
rect 43502 112338 43586 112574
rect 43822 112338 77266 112574
rect 77502 112338 77586 112574
rect 77822 112338 111266 112574
rect 111502 112338 111586 112574
rect 111822 112338 179266 112574
rect 179502 112338 179586 112574
rect 179822 112338 213266 112574
rect 213502 112338 213586 112574
rect 213822 112338 247266 112574
rect 247502 112338 247586 112574
rect 247822 112338 281266 112574
rect 281502 112338 281586 112574
rect 281822 112338 315266 112574
rect 315502 112338 315586 112574
rect 315822 112338 349266 112574
rect 349502 112338 349586 112574
rect 349822 112338 383266 112574
rect 383502 112338 383586 112574
rect 383822 112338 417266 112574
rect 417502 112338 417586 112574
rect 417822 112338 451266 112574
rect 451502 112338 451586 112574
rect 451822 112338 485266 112574
rect 485502 112338 485586 112574
rect 485822 112338 519266 112574
rect 519502 112338 519586 112574
rect 519822 112338 553266 112574
rect 553502 112338 553586 112574
rect 553822 112338 587262 112574
rect 587498 112338 587582 112574
rect 587818 112338 592650 112574
rect -8726 112306 592650 112338
rect -8726 109174 592650 109206
rect -8726 108938 -2934 109174
rect -2698 108938 -2614 109174
rect -2378 108938 5546 109174
rect 5782 108938 5866 109174
rect 6102 108938 39546 109174
rect 39782 108938 39866 109174
rect 40102 108938 73546 109174
rect 73782 108938 73866 109174
rect 74102 108938 107546 109174
rect 107782 108938 107866 109174
rect 108102 108938 135610 109174
rect 135846 108938 166330 109174
rect 166566 108938 175546 109174
rect 175782 108938 175866 109174
rect 176102 108938 209546 109174
rect 209782 108938 209866 109174
rect 210102 108938 243546 109174
rect 243782 108938 243866 109174
rect 244102 108938 277546 109174
rect 277782 108938 277866 109174
rect 278102 108938 311546 109174
rect 311782 108938 311866 109174
rect 312102 108938 345546 109174
rect 345782 108938 345866 109174
rect 346102 108938 379546 109174
rect 379782 108938 379866 109174
rect 380102 108938 413546 109174
rect 413782 108938 413866 109174
rect 414102 108938 447546 109174
rect 447782 108938 447866 109174
rect 448102 108938 481546 109174
rect 481782 108938 481866 109174
rect 482102 108938 515546 109174
rect 515782 108938 515866 109174
rect 516102 108938 549546 109174
rect 549782 108938 549866 109174
rect 550102 108938 586302 109174
rect 586538 108938 586622 109174
rect 586858 108938 592650 109174
rect -8726 108854 592650 108938
rect -8726 108618 -2934 108854
rect -2698 108618 -2614 108854
rect -2378 108618 5546 108854
rect 5782 108618 5866 108854
rect 6102 108618 39546 108854
rect 39782 108618 39866 108854
rect 40102 108618 73546 108854
rect 73782 108618 73866 108854
rect 74102 108618 107546 108854
rect 107782 108618 107866 108854
rect 108102 108618 135610 108854
rect 135846 108618 166330 108854
rect 166566 108618 175546 108854
rect 175782 108618 175866 108854
rect 176102 108618 209546 108854
rect 209782 108618 209866 108854
rect 210102 108618 243546 108854
rect 243782 108618 243866 108854
rect 244102 108618 277546 108854
rect 277782 108618 277866 108854
rect 278102 108618 311546 108854
rect 311782 108618 311866 108854
rect 312102 108618 345546 108854
rect 345782 108618 345866 108854
rect 346102 108618 379546 108854
rect 379782 108618 379866 108854
rect 380102 108618 413546 108854
rect 413782 108618 413866 108854
rect 414102 108618 447546 108854
rect 447782 108618 447866 108854
rect 448102 108618 481546 108854
rect 481782 108618 481866 108854
rect 482102 108618 515546 108854
rect 515782 108618 515866 108854
rect 516102 108618 549546 108854
rect 549782 108618 549866 108854
rect 550102 108618 586302 108854
rect 586538 108618 586622 108854
rect 586858 108618 592650 108854
rect -8726 108586 592650 108618
rect -8726 105454 592650 105486
rect -8726 105218 -1974 105454
rect -1738 105218 -1654 105454
rect -1418 105218 1826 105454
rect 2062 105218 2146 105454
rect 2382 105218 35826 105454
rect 36062 105218 36146 105454
rect 36382 105218 69826 105454
rect 70062 105218 70146 105454
rect 70382 105218 103826 105454
rect 104062 105218 104146 105454
rect 104382 105218 120250 105454
rect 120486 105218 150970 105454
rect 151206 105218 171826 105454
rect 172062 105218 172146 105454
rect 172382 105218 205826 105454
rect 206062 105218 206146 105454
rect 206382 105218 239826 105454
rect 240062 105218 240146 105454
rect 240382 105218 273826 105454
rect 274062 105218 274146 105454
rect 274382 105218 307826 105454
rect 308062 105218 308146 105454
rect 308382 105218 341826 105454
rect 342062 105218 342146 105454
rect 342382 105218 375826 105454
rect 376062 105218 376146 105454
rect 376382 105218 409826 105454
rect 410062 105218 410146 105454
rect 410382 105218 443826 105454
rect 444062 105218 444146 105454
rect 444382 105218 477826 105454
rect 478062 105218 478146 105454
rect 478382 105218 511826 105454
rect 512062 105218 512146 105454
rect 512382 105218 545826 105454
rect 546062 105218 546146 105454
rect 546382 105218 579826 105454
rect 580062 105218 580146 105454
rect 580382 105218 585342 105454
rect 585578 105218 585662 105454
rect 585898 105218 592650 105454
rect -8726 105134 592650 105218
rect -8726 104898 -1974 105134
rect -1738 104898 -1654 105134
rect -1418 104898 1826 105134
rect 2062 104898 2146 105134
rect 2382 104898 35826 105134
rect 36062 104898 36146 105134
rect 36382 104898 69826 105134
rect 70062 104898 70146 105134
rect 70382 104898 103826 105134
rect 104062 104898 104146 105134
rect 104382 104898 120250 105134
rect 120486 104898 150970 105134
rect 151206 104898 171826 105134
rect 172062 104898 172146 105134
rect 172382 104898 205826 105134
rect 206062 104898 206146 105134
rect 206382 104898 239826 105134
rect 240062 104898 240146 105134
rect 240382 104898 273826 105134
rect 274062 104898 274146 105134
rect 274382 104898 307826 105134
rect 308062 104898 308146 105134
rect 308382 104898 341826 105134
rect 342062 104898 342146 105134
rect 342382 104898 375826 105134
rect 376062 104898 376146 105134
rect 376382 104898 409826 105134
rect 410062 104898 410146 105134
rect 410382 104898 443826 105134
rect 444062 104898 444146 105134
rect 444382 104898 477826 105134
rect 478062 104898 478146 105134
rect 478382 104898 511826 105134
rect 512062 104898 512146 105134
rect 512382 104898 545826 105134
rect 546062 104898 546146 105134
rect 546382 104898 579826 105134
rect 580062 104898 580146 105134
rect 580382 104898 585342 105134
rect 585578 104898 585662 105134
rect 585898 104898 592650 105134
rect -8726 104866 592650 104898
rect -8726 97494 592650 97526
rect -8726 97258 -8694 97494
rect -8458 97258 -8374 97494
rect -8138 97258 27866 97494
rect 28102 97258 28186 97494
rect 28422 97258 61866 97494
rect 62102 97258 62186 97494
rect 62422 97258 95866 97494
rect 96102 97258 96186 97494
rect 96422 97258 197866 97494
rect 198102 97258 198186 97494
rect 198422 97258 231866 97494
rect 232102 97258 232186 97494
rect 232422 97258 265866 97494
rect 266102 97258 266186 97494
rect 266422 97258 299866 97494
rect 300102 97258 300186 97494
rect 300422 97258 333866 97494
rect 334102 97258 334186 97494
rect 334422 97258 367866 97494
rect 368102 97258 368186 97494
rect 368422 97258 401866 97494
rect 402102 97258 402186 97494
rect 402422 97258 435866 97494
rect 436102 97258 436186 97494
rect 436422 97258 469866 97494
rect 470102 97258 470186 97494
rect 470422 97258 503866 97494
rect 504102 97258 504186 97494
rect 504422 97258 537866 97494
rect 538102 97258 538186 97494
rect 538422 97258 571866 97494
rect 572102 97258 572186 97494
rect 572422 97258 592062 97494
rect 592298 97258 592382 97494
rect 592618 97258 592650 97494
rect -8726 97174 592650 97258
rect -8726 96938 -8694 97174
rect -8458 96938 -8374 97174
rect -8138 96938 27866 97174
rect 28102 96938 28186 97174
rect 28422 96938 61866 97174
rect 62102 96938 62186 97174
rect 62422 96938 95866 97174
rect 96102 96938 96186 97174
rect 96422 96938 197866 97174
rect 198102 96938 198186 97174
rect 198422 96938 231866 97174
rect 232102 96938 232186 97174
rect 232422 96938 265866 97174
rect 266102 96938 266186 97174
rect 266422 96938 299866 97174
rect 300102 96938 300186 97174
rect 300422 96938 333866 97174
rect 334102 96938 334186 97174
rect 334422 96938 367866 97174
rect 368102 96938 368186 97174
rect 368422 96938 401866 97174
rect 402102 96938 402186 97174
rect 402422 96938 435866 97174
rect 436102 96938 436186 97174
rect 436422 96938 469866 97174
rect 470102 96938 470186 97174
rect 470422 96938 503866 97174
rect 504102 96938 504186 97174
rect 504422 96938 537866 97174
rect 538102 96938 538186 97174
rect 538422 96938 571866 97174
rect 572102 96938 572186 97174
rect 572422 96938 592062 97174
rect 592298 96938 592382 97174
rect 592618 96938 592650 97174
rect -8726 96906 592650 96938
rect -8726 93774 592650 93806
rect -8726 93538 -7734 93774
rect -7498 93538 -7414 93774
rect -7178 93538 24146 93774
rect 24382 93538 24466 93774
rect 24702 93538 58146 93774
rect 58382 93538 58466 93774
rect 58702 93538 92146 93774
rect 92382 93538 92466 93774
rect 92702 93538 194146 93774
rect 194382 93538 194466 93774
rect 194702 93538 228146 93774
rect 228382 93538 228466 93774
rect 228702 93538 262146 93774
rect 262382 93538 262466 93774
rect 262702 93538 296146 93774
rect 296382 93538 296466 93774
rect 296702 93538 330146 93774
rect 330382 93538 330466 93774
rect 330702 93538 364146 93774
rect 364382 93538 364466 93774
rect 364702 93538 398146 93774
rect 398382 93538 398466 93774
rect 398702 93538 432146 93774
rect 432382 93538 432466 93774
rect 432702 93538 466146 93774
rect 466382 93538 466466 93774
rect 466702 93538 500146 93774
rect 500382 93538 500466 93774
rect 500702 93538 534146 93774
rect 534382 93538 534466 93774
rect 534702 93538 568146 93774
rect 568382 93538 568466 93774
rect 568702 93538 591102 93774
rect 591338 93538 591422 93774
rect 591658 93538 592650 93774
rect -8726 93454 592650 93538
rect -8726 93218 -7734 93454
rect -7498 93218 -7414 93454
rect -7178 93218 24146 93454
rect 24382 93218 24466 93454
rect 24702 93218 58146 93454
rect 58382 93218 58466 93454
rect 58702 93218 92146 93454
rect 92382 93218 92466 93454
rect 92702 93218 194146 93454
rect 194382 93218 194466 93454
rect 194702 93218 228146 93454
rect 228382 93218 228466 93454
rect 228702 93218 262146 93454
rect 262382 93218 262466 93454
rect 262702 93218 296146 93454
rect 296382 93218 296466 93454
rect 296702 93218 330146 93454
rect 330382 93218 330466 93454
rect 330702 93218 364146 93454
rect 364382 93218 364466 93454
rect 364702 93218 398146 93454
rect 398382 93218 398466 93454
rect 398702 93218 432146 93454
rect 432382 93218 432466 93454
rect 432702 93218 466146 93454
rect 466382 93218 466466 93454
rect 466702 93218 500146 93454
rect 500382 93218 500466 93454
rect 500702 93218 534146 93454
rect 534382 93218 534466 93454
rect 534702 93218 568146 93454
rect 568382 93218 568466 93454
rect 568702 93218 591102 93454
rect 591338 93218 591422 93454
rect 591658 93218 592650 93454
rect -8726 93186 592650 93218
rect -8726 90054 592650 90086
rect -8726 89818 -6774 90054
rect -6538 89818 -6454 90054
rect -6218 89818 20426 90054
rect 20662 89818 20746 90054
rect 20982 89818 54426 90054
rect 54662 89818 54746 90054
rect 54982 89818 88426 90054
rect 88662 89818 88746 90054
rect 88982 89818 190426 90054
rect 190662 89818 190746 90054
rect 190982 89818 224426 90054
rect 224662 89818 224746 90054
rect 224982 89818 258426 90054
rect 258662 89818 258746 90054
rect 258982 89818 292426 90054
rect 292662 89818 292746 90054
rect 292982 89818 326426 90054
rect 326662 89818 326746 90054
rect 326982 89818 360426 90054
rect 360662 89818 360746 90054
rect 360982 89818 394426 90054
rect 394662 89818 394746 90054
rect 394982 89818 428426 90054
rect 428662 89818 428746 90054
rect 428982 89818 462426 90054
rect 462662 89818 462746 90054
rect 462982 89818 496426 90054
rect 496662 89818 496746 90054
rect 496982 89818 530426 90054
rect 530662 89818 530746 90054
rect 530982 89818 564426 90054
rect 564662 89818 564746 90054
rect 564982 89818 590142 90054
rect 590378 89818 590462 90054
rect 590698 89818 592650 90054
rect -8726 89734 592650 89818
rect -8726 89498 -6774 89734
rect -6538 89498 -6454 89734
rect -6218 89498 20426 89734
rect 20662 89498 20746 89734
rect 20982 89498 54426 89734
rect 54662 89498 54746 89734
rect 54982 89498 88426 89734
rect 88662 89498 88746 89734
rect 88982 89498 190426 89734
rect 190662 89498 190746 89734
rect 190982 89498 224426 89734
rect 224662 89498 224746 89734
rect 224982 89498 258426 89734
rect 258662 89498 258746 89734
rect 258982 89498 292426 89734
rect 292662 89498 292746 89734
rect 292982 89498 326426 89734
rect 326662 89498 326746 89734
rect 326982 89498 360426 89734
rect 360662 89498 360746 89734
rect 360982 89498 394426 89734
rect 394662 89498 394746 89734
rect 394982 89498 428426 89734
rect 428662 89498 428746 89734
rect 428982 89498 462426 89734
rect 462662 89498 462746 89734
rect 462982 89498 496426 89734
rect 496662 89498 496746 89734
rect 496982 89498 530426 89734
rect 530662 89498 530746 89734
rect 530982 89498 564426 89734
rect 564662 89498 564746 89734
rect 564982 89498 590142 89734
rect 590378 89498 590462 89734
rect 590698 89498 592650 89734
rect -8726 89466 592650 89498
rect -8726 86334 592650 86366
rect -8726 86098 -5814 86334
rect -5578 86098 -5494 86334
rect -5258 86098 16706 86334
rect 16942 86098 17026 86334
rect 17262 86098 50706 86334
rect 50942 86098 51026 86334
rect 51262 86098 84706 86334
rect 84942 86098 85026 86334
rect 85262 86098 186706 86334
rect 186942 86098 187026 86334
rect 187262 86098 220706 86334
rect 220942 86098 221026 86334
rect 221262 86098 254706 86334
rect 254942 86098 255026 86334
rect 255262 86098 288706 86334
rect 288942 86098 289026 86334
rect 289262 86098 322706 86334
rect 322942 86098 323026 86334
rect 323262 86098 356706 86334
rect 356942 86098 357026 86334
rect 357262 86098 390706 86334
rect 390942 86098 391026 86334
rect 391262 86098 424706 86334
rect 424942 86098 425026 86334
rect 425262 86098 458706 86334
rect 458942 86098 459026 86334
rect 459262 86098 492706 86334
rect 492942 86098 493026 86334
rect 493262 86098 526706 86334
rect 526942 86098 527026 86334
rect 527262 86098 560706 86334
rect 560942 86098 561026 86334
rect 561262 86098 589182 86334
rect 589418 86098 589502 86334
rect 589738 86098 592650 86334
rect -8726 86014 592650 86098
rect -8726 85778 -5814 86014
rect -5578 85778 -5494 86014
rect -5258 85778 16706 86014
rect 16942 85778 17026 86014
rect 17262 85778 50706 86014
rect 50942 85778 51026 86014
rect 51262 85778 84706 86014
rect 84942 85778 85026 86014
rect 85262 85778 186706 86014
rect 186942 85778 187026 86014
rect 187262 85778 220706 86014
rect 220942 85778 221026 86014
rect 221262 85778 254706 86014
rect 254942 85778 255026 86014
rect 255262 85778 288706 86014
rect 288942 85778 289026 86014
rect 289262 85778 322706 86014
rect 322942 85778 323026 86014
rect 323262 85778 356706 86014
rect 356942 85778 357026 86014
rect 357262 85778 390706 86014
rect 390942 85778 391026 86014
rect 391262 85778 424706 86014
rect 424942 85778 425026 86014
rect 425262 85778 458706 86014
rect 458942 85778 459026 86014
rect 459262 85778 492706 86014
rect 492942 85778 493026 86014
rect 493262 85778 526706 86014
rect 526942 85778 527026 86014
rect 527262 85778 560706 86014
rect 560942 85778 561026 86014
rect 561262 85778 589182 86014
rect 589418 85778 589502 86014
rect 589738 85778 592650 86014
rect -8726 85746 592650 85778
rect -8726 82614 592650 82646
rect -8726 82378 -4854 82614
rect -4618 82378 -4534 82614
rect -4298 82378 12986 82614
rect 13222 82378 13306 82614
rect 13542 82378 46986 82614
rect 47222 82378 47306 82614
rect 47542 82378 80986 82614
rect 81222 82378 81306 82614
rect 81542 82378 114986 82614
rect 115222 82378 115306 82614
rect 115542 82378 182986 82614
rect 183222 82378 183306 82614
rect 183542 82378 216986 82614
rect 217222 82378 217306 82614
rect 217542 82378 250986 82614
rect 251222 82378 251306 82614
rect 251542 82378 284986 82614
rect 285222 82378 285306 82614
rect 285542 82378 318986 82614
rect 319222 82378 319306 82614
rect 319542 82378 352986 82614
rect 353222 82378 353306 82614
rect 353542 82378 386986 82614
rect 387222 82378 387306 82614
rect 387542 82378 420986 82614
rect 421222 82378 421306 82614
rect 421542 82378 454986 82614
rect 455222 82378 455306 82614
rect 455542 82378 488986 82614
rect 489222 82378 489306 82614
rect 489542 82378 522986 82614
rect 523222 82378 523306 82614
rect 523542 82378 556986 82614
rect 557222 82378 557306 82614
rect 557542 82378 588222 82614
rect 588458 82378 588542 82614
rect 588778 82378 592650 82614
rect -8726 82294 592650 82378
rect -8726 82058 -4854 82294
rect -4618 82058 -4534 82294
rect -4298 82058 12986 82294
rect 13222 82058 13306 82294
rect 13542 82058 46986 82294
rect 47222 82058 47306 82294
rect 47542 82058 80986 82294
rect 81222 82058 81306 82294
rect 81542 82058 114986 82294
rect 115222 82058 115306 82294
rect 115542 82058 182986 82294
rect 183222 82058 183306 82294
rect 183542 82058 216986 82294
rect 217222 82058 217306 82294
rect 217542 82058 250986 82294
rect 251222 82058 251306 82294
rect 251542 82058 284986 82294
rect 285222 82058 285306 82294
rect 285542 82058 318986 82294
rect 319222 82058 319306 82294
rect 319542 82058 352986 82294
rect 353222 82058 353306 82294
rect 353542 82058 386986 82294
rect 387222 82058 387306 82294
rect 387542 82058 420986 82294
rect 421222 82058 421306 82294
rect 421542 82058 454986 82294
rect 455222 82058 455306 82294
rect 455542 82058 488986 82294
rect 489222 82058 489306 82294
rect 489542 82058 522986 82294
rect 523222 82058 523306 82294
rect 523542 82058 556986 82294
rect 557222 82058 557306 82294
rect 557542 82058 588222 82294
rect 588458 82058 588542 82294
rect 588778 82058 592650 82294
rect -8726 82026 592650 82058
rect -8726 78894 592650 78926
rect -8726 78658 -3894 78894
rect -3658 78658 -3574 78894
rect -3338 78658 9266 78894
rect 9502 78658 9586 78894
rect 9822 78658 43266 78894
rect 43502 78658 43586 78894
rect 43822 78658 77266 78894
rect 77502 78658 77586 78894
rect 77822 78658 111266 78894
rect 111502 78658 111586 78894
rect 111822 78658 179266 78894
rect 179502 78658 179586 78894
rect 179822 78658 213266 78894
rect 213502 78658 213586 78894
rect 213822 78658 247266 78894
rect 247502 78658 247586 78894
rect 247822 78658 281266 78894
rect 281502 78658 281586 78894
rect 281822 78658 315266 78894
rect 315502 78658 315586 78894
rect 315822 78658 349266 78894
rect 349502 78658 349586 78894
rect 349822 78658 383266 78894
rect 383502 78658 383586 78894
rect 383822 78658 417266 78894
rect 417502 78658 417586 78894
rect 417822 78658 451266 78894
rect 451502 78658 451586 78894
rect 451822 78658 485266 78894
rect 485502 78658 485586 78894
rect 485822 78658 519266 78894
rect 519502 78658 519586 78894
rect 519822 78658 553266 78894
rect 553502 78658 553586 78894
rect 553822 78658 587262 78894
rect 587498 78658 587582 78894
rect 587818 78658 592650 78894
rect -8726 78574 592650 78658
rect -8726 78338 -3894 78574
rect -3658 78338 -3574 78574
rect -3338 78338 9266 78574
rect 9502 78338 9586 78574
rect 9822 78338 43266 78574
rect 43502 78338 43586 78574
rect 43822 78338 77266 78574
rect 77502 78338 77586 78574
rect 77822 78338 111266 78574
rect 111502 78338 111586 78574
rect 111822 78338 179266 78574
rect 179502 78338 179586 78574
rect 179822 78338 213266 78574
rect 213502 78338 213586 78574
rect 213822 78338 247266 78574
rect 247502 78338 247586 78574
rect 247822 78338 281266 78574
rect 281502 78338 281586 78574
rect 281822 78338 315266 78574
rect 315502 78338 315586 78574
rect 315822 78338 349266 78574
rect 349502 78338 349586 78574
rect 349822 78338 383266 78574
rect 383502 78338 383586 78574
rect 383822 78338 417266 78574
rect 417502 78338 417586 78574
rect 417822 78338 451266 78574
rect 451502 78338 451586 78574
rect 451822 78338 485266 78574
rect 485502 78338 485586 78574
rect 485822 78338 519266 78574
rect 519502 78338 519586 78574
rect 519822 78338 553266 78574
rect 553502 78338 553586 78574
rect 553822 78338 587262 78574
rect 587498 78338 587582 78574
rect 587818 78338 592650 78574
rect -8726 78306 592650 78338
rect -8726 75174 592650 75206
rect -8726 74938 -2934 75174
rect -2698 74938 -2614 75174
rect -2378 74938 5546 75174
rect 5782 74938 5866 75174
rect 6102 74938 39546 75174
rect 39782 74938 39866 75174
rect 40102 74938 73546 75174
rect 73782 74938 73866 75174
rect 74102 74938 107546 75174
rect 107782 74938 107866 75174
rect 108102 74938 175546 75174
rect 175782 74938 175866 75174
rect 176102 74938 209546 75174
rect 209782 74938 209866 75174
rect 210102 74938 243546 75174
rect 243782 74938 243866 75174
rect 244102 74938 277546 75174
rect 277782 74938 277866 75174
rect 278102 74938 311546 75174
rect 311782 74938 311866 75174
rect 312102 74938 345546 75174
rect 345782 74938 345866 75174
rect 346102 74938 379546 75174
rect 379782 74938 379866 75174
rect 380102 74938 413546 75174
rect 413782 74938 413866 75174
rect 414102 74938 447546 75174
rect 447782 74938 447866 75174
rect 448102 74938 481546 75174
rect 481782 74938 481866 75174
rect 482102 74938 515546 75174
rect 515782 74938 515866 75174
rect 516102 74938 549546 75174
rect 549782 74938 549866 75174
rect 550102 74938 586302 75174
rect 586538 74938 586622 75174
rect 586858 74938 592650 75174
rect -8726 74854 592650 74938
rect -8726 74618 -2934 74854
rect -2698 74618 -2614 74854
rect -2378 74618 5546 74854
rect 5782 74618 5866 74854
rect 6102 74618 39546 74854
rect 39782 74618 39866 74854
rect 40102 74618 73546 74854
rect 73782 74618 73866 74854
rect 74102 74618 107546 74854
rect 107782 74618 107866 74854
rect 108102 74618 175546 74854
rect 175782 74618 175866 74854
rect 176102 74618 209546 74854
rect 209782 74618 209866 74854
rect 210102 74618 243546 74854
rect 243782 74618 243866 74854
rect 244102 74618 277546 74854
rect 277782 74618 277866 74854
rect 278102 74618 311546 74854
rect 311782 74618 311866 74854
rect 312102 74618 345546 74854
rect 345782 74618 345866 74854
rect 346102 74618 379546 74854
rect 379782 74618 379866 74854
rect 380102 74618 413546 74854
rect 413782 74618 413866 74854
rect 414102 74618 447546 74854
rect 447782 74618 447866 74854
rect 448102 74618 481546 74854
rect 481782 74618 481866 74854
rect 482102 74618 515546 74854
rect 515782 74618 515866 74854
rect 516102 74618 549546 74854
rect 549782 74618 549866 74854
rect 550102 74618 586302 74854
rect 586538 74618 586622 74854
rect 586858 74618 592650 74854
rect -8726 74586 592650 74618
rect -8726 71454 592650 71486
rect -8726 71218 -1974 71454
rect -1738 71218 -1654 71454
rect -1418 71218 1826 71454
rect 2062 71218 2146 71454
rect 2382 71218 35826 71454
rect 36062 71218 36146 71454
rect 36382 71218 69826 71454
rect 70062 71218 70146 71454
rect 70382 71218 103826 71454
rect 104062 71218 104146 71454
rect 104382 71218 137826 71454
rect 138062 71218 138146 71454
rect 138382 71218 171826 71454
rect 172062 71218 172146 71454
rect 172382 71218 205826 71454
rect 206062 71218 206146 71454
rect 206382 71218 239826 71454
rect 240062 71218 240146 71454
rect 240382 71218 273826 71454
rect 274062 71218 274146 71454
rect 274382 71218 307826 71454
rect 308062 71218 308146 71454
rect 308382 71218 341826 71454
rect 342062 71218 342146 71454
rect 342382 71218 375826 71454
rect 376062 71218 376146 71454
rect 376382 71218 409826 71454
rect 410062 71218 410146 71454
rect 410382 71218 443826 71454
rect 444062 71218 444146 71454
rect 444382 71218 477826 71454
rect 478062 71218 478146 71454
rect 478382 71218 511826 71454
rect 512062 71218 512146 71454
rect 512382 71218 545826 71454
rect 546062 71218 546146 71454
rect 546382 71218 579826 71454
rect 580062 71218 580146 71454
rect 580382 71218 585342 71454
rect 585578 71218 585662 71454
rect 585898 71218 592650 71454
rect -8726 71134 592650 71218
rect -8726 70898 -1974 71134
rect -1738 70898 -1654 71134
rect -1418 70898 1826 71134
rect 2062 70898 2146 71134
rect 2382 70898 35826 71134
rect 36062 70898 36146 71134
rect 36382 70898 69826 71134
rect 70062 70898 70146 71134
rect 70382 70898 103826 71134
rect 104062 70898 104146 71134
rect 104382 70898 137826 71134
rect 138062 70898 138146 71134
rect 138382 70898 171826 71134
rect 172062 70898 172146 71134
rect 172382 70898 205826 71134
rect 206062 70898 206146 71134
rect 206382 70898 239826 71134
rect 240062 70898 240146 71134
rect 240382 70898 273826 71134
rect 274062 70898 274146 71134
rect 274382 70898 307826 71134
rect 308062 70898 308146 71134
rect 308382 70898 341826 71134
rect 342062 70898 342146 71134
rect 342382 70898 375826 71134
rect 376062 70898 376146 71134
rect 376382 70898 409826 71134
rect 410062 70898 410146 71134
rect 410382 70898 443826 71134
rect 444062 70898 444146 71134
rect 444382 70898 477826 71134
rect 478062 70898 478146 71134
rect 478382 70898 511826 71134
rect 512062 70898 512146 71134
rect 512382 70898 545826 71134
rect 546062 70898 546146 71134
rect 546382 70898 579826 71134
rect 580062 70898 580146 71134
rect 580382 70898 585342 71134
rect 585578 70898 585662 71134
rect 585898 70898 592650 71134
rect -8726 70866 592650 70898
rect -8726 63494 592650 63526
rect -8726 63258 -8694 63494
rect -8458 63258 -8374 63494
rect -8138 63258 27866 63494
rect 28102 63258 28186 63494
rect 28422 63258 61866 63494
rect 62102 63258 62186 63494
rect 62422 63258 95866 63494
rect 96102 63258 96186 63494
rect 96422 63258 129866 63494
rect 130102 63258 130186 63494
rect 130422 63258 163866 63494
rect 164102 63258 164186 63494
rect 164422 63258 197866 63494
rect 198102 63258 198186 63494
rect 198422 63258 231866 63494
rect 232102 63258 232186 63494
rect 232422 63258 265866 63494
rect 266102 63258 266186 63494
rect 266422 63258 299866 63494
rect 300102 63258 300186 63494
rect 300422 63258 333866 63494
rect 334102 63258 334186 63494
rect 334422 63258 367866 63494
rect 368102 63258 368186 63494
rect 368422 63258 401866 63494
rect 402102 63258 402186 63494
rect 402422 63258 435866 63494
rect 436102 63258 436186 63494
rect 436422 63258 469866 63494
rect 470102 63258 470186 63494
rect 470422 63258 503866 63494
rect 504102 63258 504186 63494
rect 504422 63258 537866 63494
rect 538102 63258 538186 63494
rect 538422 63258 571866 63494
rect 572102 63258 572186 63494
rect 572422 63258 592062 63494
rect 592298 63258 592382 63494
rect 592618 63258 592650 63494
rect -8726 63174 592650 63258
rect -8726 62938 -8694 63174
rect -8458 62938 -8374 63174
rect -8138 62938 27866 63174
rect 28102 62938 28186 63174
rect 28422 62938 61866 63174
rect 62102 62938 62186 63174
rect 62422 62938 95866 63174
rect 96102 62938 96186 63174
rect 96422 62938 129866 63174
rect 130102 62938 130186 63174
rect 130422 62938 163866 63174
rect 164102 62938 164186 63174
rect 164422 62938 197866 63174
rect 198102 62938 198186 63174
rect 198422 62938 231866 63174
rect 232102 62938 232186 63174
rect 232422 62938 265866 63174
rect 266102 62938 266186 63174
rect 266422 62938 299866 63174
rect 300102 62938 300186 63174
rect 300422 62938 333866 63174
rect 334102 62938 334186 63174
rect 334422 62938 367866 63174
rect 368102 62938 368186 63174
rect 368422 62938 401866 63174
rect 402102 62938 402186 63174
rect 402422 62938 435866 63174
rect 436102 62938 436186 63174
rect 436422 62938 469866 63174
rect 470102 62938 470186 63174
rect 470422 62938 503866 63174
rect 504102 62938 504186 63174
rect 504422 62938 537866 63174
rect 538102 62938 538186 63174
rect 538422 62938 571866 63174
rect 572102 62938 572186 63174
rect 572422 62938 592062 63174
rect 592298 62938 592382 63174
rect 592618 62938 592650 63174
rect -8726 62906 592650 62938
rect -8726 59774 592650 59806
rect -8726 59538 -7734 59774
rect -7498 59538 -7414 59774
rect -7178 59538 24146 59774
rect 24382 59538 24466 59774
rect 24702 59538 58146 59774
rect 58382 59538 58466 59774
rect 58702 59538 92146 59774
rect 92382 59538 92466 59774
rect 92702 59538 126146 59774
rect 126382 59538 126466 59774
rect 126702 59538 160146 59774
rect 160382 59538 160466 59774
rect 160702 59538 194146 59774
rect 194382 59538 194466 59774
rect 194702 59538 228146 59774
rect 228382 59538 228466 59774
rect 228702 59538 262146 59774
rect 262382 59538 262466 59774
rect 262702 59538 296146 59774
rect 296382 59538 296466 59774
rect 296702 59538 330146 59774
rect 330382 59538 330466 59774
rect 330702 59538 364146 59774
rect 364382 59538 364466 59774
rect 364702 59538 398146 59774
rect 398382 59538 398466 59774
rect 398702 59538 432146 59774
rect 432382 59538 432466 59774
rect 432702 59538 466146 59774
rect 466382 59538 466466 59774
rect 466702 59538 500146 59774
rect 500382 59538 500466 59774
rect 500702 59538 534146 59774
rect 534382 59538 534466 59774
rect 534702 59538 568146 59774
rect 568382 59538 568466 59774
rect 568702 59538 591102 59774
rect 591338 59538 591422 59774
rect 591658 59538 592650 59774
rect -8726 59454 592650 59538
rect -8726 59218 -7734 59454
rect -7498 59218 -7414 59454
rect -7178 59218 24146 59454
rect 24382 59218 24466 59454
rect 24702 59218 58146 59454
rect 58382 59218 58466 59454
rect 58702 59218 92146 59454
rect 92382 59218 92466 59454
rect 92702 59218 126146 59454
rect 126382 59218 126466 59454
rect 126702 59218 160146 59454
rect 160382 59218 160466 59454
rect 160702 59218 194146 59454
rect 194382 59218 194466 59454
rect 194702 59218 228146 59454
rect 228382 59218 228466 59454
rect 228702 59218 262146 59454
rect 262382 59218 262466 59454
rect 262702 59218 296146 59454
rect 296382 59218 296466 59454
rect 296702 59218 330146 59454
rect 330382 59218 330466 59454
rect 330702 59218 364146 59454
rect 364382 59218 364466 59454
rect 364702 59218 398146 59454
rect 398382 59218 398466 59454
rect 398702 59218 432146 59454
rect 432382 59218 432466 59454
rect 432702 59218 466146 59454
rect 466382 59218 466466 59454
rect 466702 59218 500146 59454
rect 500382 59218 500466 59454
rect 500702 59218 534146 59454
rect 534382 59218 534466 59454
rect 534702 59218 568146 59454
rect 568382 59218 568466 59454
rect 568702 59218 591102 59454
rect 591338 59218 591422 59454
rect 591658 59218 592650 59454
rect -8726 59186 592650 59218
rect -8726 56054 592650 56086
rect -8726 55818 -6774 56054
rect -6538 55818 -6454 56054
rect -6218 55818 20426 56054
rect 20662 55818 20746 56054
rect 20982 55818 54426 56054
rect 54662 55818 54746 56054
rect 54982 55818 88426 56054
rect 88662 55818 88746 56054
rect 88982 55818 122426 56054
rect 122662 55818 122746 56054
rect 122982 55818 156426 56054
rect 156662 55818 156746 56054
rect 156982 55818 190426 56054
rect 190662 55818 190746 56054
rect 190982 55818 224426 56054
rect 224662 55818 224746 56054
rect 224982 55818 258426 56054
rect 258662 55818 258746 56054
rect 258982 55818 292426 56054
rect 292662 55818 292746 56054
rect 292982 55818 326426 56054
rect 326662 55818 326746 56054
rect 326982 55818 360426 56054
rect 360662 55818 360746 56054
rect 360982 55818 394426 56054
rect 394662 55818 394746 56054
rect 394982 55818 428426 56054
rect 428662 55818 428746 56054
rect 428982 55818 462426 56054
rect 462662 55818 462746 56054
rect 462982 55818 496426 56054
rect 496662 55818 496746 56054
rect 496982 55818 530426 56054
rect 530662 55818 530746 56054
rect 530982 55818 564426 56054
rect 564662 55818 564746 56054
rect 564982 55818 590142 56054
rect 590378 55818 590462 56054
rect 590698 55818 592650 56054
rect -8726 55734 592650 55818
rect -8726 55498 -6774 55734
rect -6538 55498 -6454 55734
rect -6218 55498 20426 55734
rect 20662 55498 20746 55734
rect 20982 55498 54426 55734
rect 54662 55498 54746 55734
rect 54982 55498 88426 55734
rect 88662 55498 88746 55734
rect 88982 55498 122426 55734
rect 122662 55498 122746 55734
rect 122982 55498 156426 55734
rect 156662 55498 156746 55734
rect 156982 55498 190426 55734
rect 190662 55498 190746 55734
rect 190982 55498 224426 55734
rect 224662 55498 224746 55734
rect 224982 55498 258426 55734
rect 258662 55498 258746 55734
rect 258982 55498 292426 55734
rect 292662 55498 292746 55734
rect 292982 55498 326426 55734
rect 326662 55498 326746 55734
rect 326982 55498 360426 55734
rect 360662 55498 360746 55734
rect 360982 55498 394426 55734
rect 394662 55498 394746 55734
rect 394982 55498 428426 55734
rect 428662 55498 428746 55734
rect 428982 55498 462426 55734
rect 462662 55498 462746 55734
rect 462982 55498 496426 55734
rect 496662 55498 496746 55734
rect 496982 55498 530426 55734
rect 530662 55498 530746 55734
rect 530982 55498 564426 55734
rect 564662 55498 564746 55734
rect 564982 55498 590142 55734
rect 590378 55498 590462 55734
rect 590698 55498 592650 55734
rect -8726 55466 592650 55498
rect -8726 52334 592650 52366
rect -8726 52098 -5814 52334
rect -5578 52098 -5494 52334
rect -5258 52098 16706 52334
rect 16942 52098 17026 52334
rect 17262 52098 50706 52334
rect 50942 52098 51026 52334
rect 51262 52098 84706 52334
rect 84942 52098 85026 52334
rect 85262 52098 118706 52334
rect 118942 52098 119026 52334
rect 119262 52098 152706 52334
rect 152942 52098 153026 52334
rect 153262 52098 186706 52334
rect 186942 52098 187026 52334
rect 187262 52098 220706 52334
rect 220942 52098 221026 52334
rect 221262 52098 254706 52334
rect 254942 52098 255026 52334
rect 255262 52098 288706 52334
rect 288942 52098 289026 52334
rect 289262 52098 322706 52334
rect 322942 52098 323026 52334
rect 323262 52098 356706 52334
rect 356942 52098 357026 52334
rect 357262 52098 390706 52334
rect 390942 52098 391026 52334
rect 391262 52098 424706 52334
rect 424942 52098 425026 52334
rect 425262 52098 458706 52334
rect 458942 52098 459026 52334
rect 459262 52098 492706 52334
rect 492942 52098 493026 52334
rect 493262 52098 526706 52334
rect 526942 52098 527026 52334
rect 527262 52098 560706 52334
rect 560942 52098 561026 52334
rect 561262 52098 589182 52334
rect 589418 52098 589502 52334
rect 589738 52098 592650 52334
rect -8726 52014 592650 52098
rect -8726 51778 -5814 52014
rect -5578 51778 -5494 52014
rect -5258 51778 16706 52014
rect 16942 51778 17026 52014
rect 17262 51778 50706 52014
rect 50942 51778 51026 52014
rect 51262 51778 84706 52014
rect 84942 51778 85026 52014
rect 85262 51778 118706 52014
rect 118942 51778 119026 52014
rect 119262 51778 152706 52014
rect 152942 51778 153026 52014
rect 153262 51778 186706 52014
rect 186942 51778 187026 52014
rect 187262 51778 220706 52014
rect 220942 51778 221026 52014
rect 221262 51778 254706 52014
rect 254942 51778 255026 52014
rect 255262 51778 288706 52014
rect 288942 51778 289026 52014
rect 289262 51778 322706 52014
rect 322942 51778 323026 52014
rect 323262 51778 356706 52014
rect 356942 51778 357026 52014
rect 357262 51778 390706 52014
rect 390942 51778 391026 52014
rect 391262 51778 424706 52014
rect 424942 51778 425026 52014
rect 425262 51778 458706 52014
rect 458942 51778 459026 52014
rect 459262 51778 492706 52014
rect 492942 51778 493026 52014
rect 493262 51778 526706 52014
rect 526942 51778 527026 52014
rect 527262 51778 560706 52014
rect 560942 51778 561026 52014
rect 561262 51778 589182 52014
rect 589418 51778 589502 52014
rect 589738 51778 592650 52014
rect -8726 51746 592650 51778
rect -8726 48614 592650 48646
rect -8726 48378 -4854 48614
rect -4618 48378 -4534 48614
rect -4298 48378 12986 48614
rect 13222 48378 13306 48614
rect 13542 48378 46986 48614
rect 47222 48378 47306 48614
rect 47542 48378 80986 48614
rect 81222 48378 81306 48614
rect 81542 48378 114986 48614
rect 115222 48378 115306 48614
rect 115542 48378 148986 48614
rect 149222 48378 149306 48614
rect 149542 48378 182986 48614
rect 183222 48378 183306 48614
rect 183542 48378 216986 48614
rect 217222 48378 217306 48614
rect 217542 48378 250986 48614
rect 251222 48378 251306 48614
rect 251542 48378 284986 48614
rect 285222 48378 285306 48614
rect 285542 48378 318986 48614
rect 319222 48378 319306 48614
rect 319542 48378 352986 48614
rect 353222 48378 353306 48614
rect 353542 48378 386986 48614
rect 387222 48378 387306 48614
rect 387542 48378 420986 48614
rect 421222 48378 421306 48614
rect 421542 48378 454986 48614
rect 455222 48378 455306 48614
rect 455542 48378 488986 48614
rect 489222 48378 489306 48614
rect 489542 48378 522986 48614
rect 523222 48378 523306 48614
rect 523542 48378 556986 48614
rect 557222 48378 557306 48614
rect 557542 48378 588222 48614
rect 588458 48378 588542 48614
rect 588778 48378 592650 48614
rect -8726 48294 592650 48378
rect -8726 48058 -4854 48294
rect -4618 48058 -4534 48294
rect -4298 48058 12986 48294
rect 13222 48058 13306 48294
rect 13542 48058 46986 48294
rect 47222 48058 47306 48294
rect 47542 48058 80986 48294
rect 81222 48058 81306 48294
rect 81542 48058 114986 48294
rect 115222 48058 115306 48294
rect 115542 48058 148986 48294
rect 149222 48058 149306 48294
rect 149542 48058 182986 48294
rect 183222 48058 183306 48294
rect 183542 48058 216986 48294
rect 217222 48058 217306 48294
rect 217542 48058 250986 48294
rect 251222 48058 251306 48294
rect 251542 48058 284986 48294
rect 285222 48058 285306 48294
rect 285542 48058 318986 48294
rect 319222 48058 319306 48294
rect 319542 48058 352986 48294
rect 353222 48058 353306 48294
rect 353542 48058 386986 48294
rect 387222 48058 387306 48294
rect 387542 48058 420986 48294
rect 421222 48058 421306 48294
rect 421542 48058 454986 48294
rect 455222 48058 455306 48294
rect 455542 48058 488986 48294
rect 489222 48058 489306 48294
rect 489542 48058 522986 48294
rect 523222 48058 523306 48294
rect 523542 48058 556986 48294
rect 557222 48058 557306 48294
rect 557542 48058 588222 48294
rect 588458 48058 588542 48294
rect 588778 48058 592650 48294
rect -8726 48026 592650 48058
rect -8726 44894 592650 44926
rect -8726 44658 -3894 44894
rect -3658 44658 -3574 44894
rect -3338 44658 9266 44894
rect 9502 44658 9586 44894
rect 9822 44658 43266 44894
rect 43502 44658 43586 44894
rect 43822 44658 77266 44894
rect 77502 44658 77586 44894
rect 77822 44658 111266 44894
rect 111502 44658 111586 44894
rect 111822 44658 145266 44894
rect 145502 44658 145586 44894
rect 145822 44658 179266 44894
rect 179502 44658 179586 44894
rect 179822 44658 213266 44894
rect 213502 44658 213586 44894
rect 213822 44658 247266 44894
rect 247502 44658 247586 44894
rect 247822 44658 281266 44894
rect 281502 44658 281586 44894
rect 281822 44658 315266 44894
rect 315502 44658 315586 44894
rect 315822 44658 349266 44894
rect 349502 44658 349586 44894
rect 349822 44658 383266 44894
rect 383502 44658 383586 44894
rect 383822 44658 417266 44894
rect 417502 44658 417586 44894
rect 417822 44658 451266 44894
rect 451502 44658 451586 44894
rect 451822 44658 485266 44894
rect 485502 44658 485586 44894
rect 485822 44658 519266 44894
rect 519502 44658 519586 44894
rect 519822 44658 553266 44894
rect 553502 44658 553586 44894
rect 553822 44658 587262 44894
rect 587498 44658 587582 44894
rect 587818 44658 592650 44894
rect -8726 44574 592650 44658
rect -8726 44338 -3894 44574
rect -3658 44338 -3574 44574
rect -3338 44338 9266 44574
rect 9502 44338 9586 44574
rect 9822 44338 43266 44574
rect 43502 44338 43586 44574
rect 43822 44338 77266 44574
rect 77502 44338 77586 44574
rect 77822 44338 111266 44574
rect 111502 44338 111586 44574
rect 111822 44338 145266 44574
rect 145502 44338 145586 44574
rect 145822 44338 179266 44574
rect 179502 44338 179586 44574
rect 179822 44338 213266 44574
rect 213502 44338 213586 44574
rect 213822 44338 247266 44574
rect 247502 44338 247586 44574
rect 247822 44338 281266 44574
rect 281502 44338 281586 44574
rect 281822 44338 315266 44574
rect 315502 44338 315586 44574
rect 315822 44338 349266 44574
rect 349502 44338 349586 44574
rect 349822 44338 383266 44574
rect 383502 44338 383586 44574
rect 383822 44338 417266 44574
rect 417502 44338 417586 44574
rect 417822 44338 451266 44574
rect 451502 44338 451586 44574
rect 451822 44338 485266 44574
rect 485502 44338 485586 44574
rect 485822 44338 519266 44574
rect 519502 44338 519586 44574
rect 519822 44338 553266 44574
rect 553502 44338 553586 44574
rect 553822 44338 587262 44574
rect 587498 44338 587582 44574
rect 587818 44338 592650 44574
rect -8726 44306 592650 44338
rect -8726 41174 592650 41206
rect -8726 40938 -2934 41174
rect -2698 40938 -2614 41174
rect -2378 40938 5546 41174
rect 5782 40938 5866 41174
rect 6102 40938 39546 41174
rect 39782 40938 39866 41174
rect 40102 40938 73546 41174
rect 73782 40938 73866 41174
rect 74102 40938 107546 41174
rect 107782 40938 107866 41174
rect 108102 40938 141546 41174
rect 141782 40938 141866 41174
rect 142102 40938 175546 41174
rect 175782 40938 175866 41174
rect 176102 40938 209546 41174
rect 209782 40938 209866 41174
rect 210102 40938 243546 41174
rect 243782 40938 243866 41174
rect 244102 40938 277546 41174
rect 277782 40938 277866 41174
rect 278102 40938 311546 41174
rect 311782 40938 311866 41174
rect 312102 40938 345546 41174
rect 345782 40938 345866 41174
rect 346102 40938 379546 41174
rect 379782 40938 379866 41174
rect 380102 40938 413546 41174
rect 413782 40938 413866 41174
rect 414102 40938 447546 41174
rect 447782 40938 447866 41174
rect 448102 40938 481546 41174
rect 481782 40938 481866 41174
rect 482102 40938 515546 41174
rect 515782 40938 515866 41174
rect 516102 40938 549546 41174
rect 549782 40938 549866 41174
rect 550102 40938 586302 41174
rect 586538 40938 586622 41174
rect 586858 40938 592650 41174
rect -8726 40854 592650 40938
rect -8726 40618 -2934 40854
rect -2698 40618 -2614 40854
rect -2378 40618 5546 40854
rect 5782 40618 5866 40854
rect 6102 40618 39546 40854
rect 39782 40618 39866 40854
rect 40102 40618 73546 40854
rect 73782 40618 73866 40854
rect 74102 40618 107546 40854
rect 107782 40618 107866 40854
rect 108102 40618 141546 40854
rect 141782 40618 141866 40854
rect 142102 40618 175546 40854
rect 175782 40618 175866 40854
rect 176102 40618 209546 40854
rect 209782 40618 209866 40854
rect 210102 40618 243546 40854
rect 243782 40618 243866 40854
rect 244102 40618 277546 40854
rect 277782 40618 277866 40854
rect 278102 40618 311546 40854
rect 311782 40618 311866 40854
rect 312102 40618 345546 40854
rect 345782 40618 345866 40854
rect 346102 40618 379546 40854
rect 379782 40618 379866 40854
rect 380102 40618 413546 40854
rect 413782 40618 413866 40854
rect 414102 40618 447546 40854
rect 447782 40618 447866 40854
rect 448102 40618 481546 40854
rect 481782 40618 481866 40854
rect 482102 40618 515546 40854
rect 515782 40618 515866 40854
rect 516102 40618 549546 40854
rect 549782 40618 549866 40854
rect 550102 40618 586302 40854
rect 586538 40618 586622 40854
rect 586858 40618 592650 40854
rect -8726 40586 592650 40618
rect -8726 37454 592650 37486
rect -8726 37218 -1974 37454
rect -1738 37218 -1654 37454
rect -1418 37218 1826 37454
rect 2062 37218 2146 37454
rect 2382 37218 35826 37454
rect 36062 37218 36146 37454
rect 36382 37218 69826 37454
rect 70062 37218 70146 37454
rect 70382 37218 103826 37454
rect 104062 37218 104146 37454
rect 104382 37218 137826 37454
rect 138062 37218 138146 37454
rect 138382 37218 171826 37454
rect 172062 37218 172146 37454
rect 172382 37218 205826 37454
rect 206062 37218 206146 37454
rect 206382 37218 239826 37454
rect 240062 37218 240146 37454
rect 240382 37218 273826 37454
rect 274062 37218 274146 37454
rect 274382 37218 307826 37454
rect 308062 37218 308146 37454
rect 308382 37218 341826 37454
rect 342062 37218 342146 37454
rect 342382 37218 375826 37454
rect 376062 37218 376146 37454
rect 376382 37218 409826 37454
rect 410062 37218 410146 37454
rect 410382 37218 443826 37454
rect 444062 37218 444146 37454
rect 444382 37218 477826 37454
rect 478062 37218 478146 37454
rect 478382 37218 511826 37454
rect 512062 37218 512146 37454
rect 512382 37218 545826 37454
rect 546062 37218 546146 37454
rect 546382 37218 579826 37454
rect 580062 37218 580146 37454
rect 580382 37218 585342 37454
rect 585578 37218 585662 37454
rect 585898 37218 592650 37454
rect -8726 37134 592650 37218
rect -8726 36898 -1974 37134
rect -1738 36898 -1654 37134
rect -1418 36898 1826 37134
rect 2062 36898 2146 37134
rect 2382 36898 35826 37134
rect 36062 36898 36146 37134
rect 36382 36898 69826 37134
rect 70062 36898 70146 37134
rect 70382 36898 103826 37134
rect 104062 36898 104146 37134
rect 104382 36898 137826 37134
rect 138062 36898 138146 37134
rect 138382 36898 171826 37134
rect 172062 36898 172146 37134
rect 172382 36898 205826 37134
rect 206062 36898 206146 37134
rect 206382 36898 239826 37134
rect 240062 36898 240146 37134
rect 240382 36898 273826 37134
rect 274062 36898 274146 37134
rect 274382 36898 307826 37134
rect 308062 36898 308146 37134
rect 308382 36898 341826 37134
rect 342062 36898 342146 37134
rect 342382 36898 375826 37134
rect 376062 36898 376146 37134
rect 376382 36898 409826 37134
rect 410062 36898 410146 37134
rect 410382 36898 443826 37134
rect 444062 36898 444146 37134
rect 444382 36898 477826 37134
rect 478062 36898 478146 37134
rect 478382 36898 511826 37134
rect 512062 36898 512146 37134
rect 512382 36898 545826 37134
rect 546062 36898 546146 37134
rect 546382 36898 579826 37134
rect 580062 36898 580146 37134
rect 580382 36898 585342 37134
rect 585578 36898 585662 37134
rect 585898 36898 592650 37134
rect -8726 36866 592650 36898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 61866 29494
rect 62102 29258 62186 29494
rect 62422 29258 95866 29494
rect 96102 29258 96186 29494
rect 96422 29258 129866 29494
rect 130102 29258 130186 29494
rect 130422 29258 163866 29494
rect 164102 29258 164186 29494
rect 164422 29258 197866 29494
rect 198102 29258 198186 29494
rect 198422 29258 231866 29494
rect 232102 29258 232186 29494
rect 232422 29258 265866 29494
rect 266102 29258 266186 29494
rect 266422 29258 299866 29494
rect 300102 29258 300186 29494
rect 300422 29258 333866 29494
rect 334102 29258 334186 29494
rect 334422 29258 367866 29494
rect 368102 29258 368186 29494
rect 368422 29258 401866 29494
rect 402102 29258 402186 29494
rect 402422 29258 435866 29494
rect 436102 29258 436186 29494
rect 436422 29258 469866 29494
rect 470102 29258 470186 29494
rect 470422 29258 503866 29494
rect 504102 29258 504186 29494
rect 504422 29258 537866 29494
rect 538102 29258 538186 29494
rect 538422 29258 571866 29494
rect 572102 29258 572186 29494
rect 572422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 61866 29174
rect 62102 28938 62186 29174
rect 62422 28938 95866 29174
rect 96102 28938 96186 29174
rect 96422 28938 129866 29174
rect 130102 28938 130186 29174
rect 130422 28938 163866 29174
rect 164102 28938 164186 29174
rect 164422 28938 197866 29174
rect 198102 28938 198186 29174
rect 198422 28938 231866 29174
rect 232102 28938 232186 29174
rect 232422 28938 265866 29174
rect 266102 28938 266186 29174
rect 266422 28938 299866 29174
rect 300102 28938 300186 29174
rect 300422 28938 333866 29174
rect 334102 28938 334186 29174
rect 334422 28938 367866 29174
rect 368102 28938 368186 29174
rect 368422 28938 401866 29174
rect 402102 28938 402186 29174
rect 402422 28938 435866 29174
rect 436102 28938 436186 29174
rect 436422 28938 469866 29174
rect 470102 28938 470186 29174
rect 470422 28938 503866 29174
rect 504102 28938 504186 29174
rect 504422 28938 537866 29174
rect 538102 28938 538186 29174
rect 538422 28938 571866 29174
rect 572102 28938 572186 29174
rect 572422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 58146 25774
rect 58382 25538 58466 25774
rect 58702 25538 92146 25774
rect 92382 25538 92466 25774
rect 92702 25538 126146 25774
rect 126382 25538 126466 25774
rect 126702 25538 160146 25774
rect 160382 25538 160466 25774
rect 160702 25538 194146 25774
rect 194382 25538 194466 25774
rect 194702 25538 228146 25774
rect 228382 25538 228466 25774
rect 228702 25538 262146 25774
rect 262382 25538 262466 25774
rect 262702 25538 296146 25774
rect 296382 25538 296466 25774
rect 296702 25538 330146 25774
rect 330382 25538 330466 25774
rect 330702 25538 364146 25774
rect 364382 25538 364466 25774
rect 364702 25538 398146 25774
rect 398382 25538 398466 25774
rect 398702 25538 432146 25774
rect 432382 25538 432466 25774
rect 432702 25538 466146 25774
rect 466382 25538 466466 25774
rect 466702 25538 500146 25774
rect 500382 25538 500466 25774
rect 500702 25538 534146 25774
rect 534382 25538 534466 25774
rect 534702 25538 568146 25774
rect 568382 25538 568466 25774
rect 568702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 58146 25454
rect 58382 25218 58466 25454
rect 58702 25218 92146 25454
rect 92382 25218 92466 25454
rect 92702 25218 126146 25454
rect 126382 25218 126466 25454
rect 126702 25218 160146 25454
rect 160382 25218 160466 25454
rect 160702 25218 194146 25454
rect 194382 25218 194466 25454
rect 194702 25218 228146 25454
rect 228382 25218 228466 25454
rect 228702 25218 262146 25454
rect 262382 25218 262466 25454
rect 262702 25218 296146 25454
rect 296382 25218 296466 25454
rect 296702 25218 330146 25454
rect 330382 25218 330466 25454
rect 330702 25218 364146 25454
rect 364382 25218 364466 25454
rect 364702 25218 398146 25454
rect 398382 25218 398466 25454
rect 398702 25218 432146 25454
rect 432382 25218 432466 25454
rect 432702 25218 466146 25454
rect 466382 25218 466466 25454
rect 466702 25218 500146 25454
rect 500382 25218 500466 25454
rect 500702 25218 534146 25454
rect 534382 25218 534466 25454
rect 534702 25218 568146 25454
rect 568382 25218 568466 25454
rect 568702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 54426 22054
rect 54662 21818 54746 22054
rect 54982 21818 88426 22054
rect 88662 21818 88746 22054
rect 88982 21818 122426 22054
rect 122662 21818 122746 22054
rect 122982 21818 156426 22054
rect 156662 21818 156746 22054
rect 156982 21818 190426 22054
rect 190662 21818 190746 22054
rect 190982 21818 224426 22054
rect 224662 21818 224746 22054
rect 224982 21818 258426 22054
rect 258662 21818 258746 22054
rect 258982 21818 292426 22054
rect 292662 21818 292746 22054
rect 292982 21818 326426 22054
rect 326662 21818 326746 22054
rect 326982 21818 360426 22054
rect 360662 21818 360746 22054
rect 360982 21818 394426 22054
rect 394662 21818 394746 22054
rect 394982 21818 428426 22054
rect 428662 21818 428746 22054
rect 428982 21818 462426 22054
rect 462662 21818 462746 22054
rect 462982 21818 496426 22054
rect 496662 21818 496746 22054
rect 496982 21818 530426 22054
rect 530662 21818 530746 22054
rect 530982 21818 564426 22054
rect 564662 21818 564746 22054
rect 564982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 54426 21734
rect 54662 21498 54746 21734
rect 54982 21498 88426 21734
rect 88662 21498 88746 21734
rect 88982 21498 122426 21734
rect 122662 21498 122746 21734
rect 122982 21498 156426 21734
rect 156662 21498 156746 21734
rect 156982 21498 190426 21734
rect 190662 21498 190746 21734
rect 190982 21498 224426 21734
rect 224662 21498 224746 21734
rect 224982 21498 258426 21734
rect 258662 21498 258746 21734
rect 258982 21498 292426 21734
rect 292662 21498 292746 21734
rect 292982 21498 326426 21734
rect 326662 21498 326746 21734
rect 326982 21498 360426 21734
rect 360662 21498 360746 21734
rect 360982 21498 394426 21734
rect 394662 21498 394746 21734
rect 394982 21498 428426 21734
rect 428662 21498 428746 21734
rect 428982 21498 462426 21734
rect 462662 21498 462746 21734
rect 462982 21498 496426 21734
rect 496662 21498 496746 21734
rect 496982 21498 530426 21734
rect 530662 21498 530746 21734
rect 530982 21498 564426 21734
rect 564662 21498 564746 21734
rect 564982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 50706 18334
rect 50942 18098 51026 18334
rect 51262 18098 84706 18334
rect 84942 18098 85026 18334
rect 85262 18098 118706 18334
rect 118942 18098 119026 18334
rect 119262 18098 152706 18334
rect 152942 18098 153026 18334
rect 153262 18098 186706 18334
rect 186942 18098 187026 18334
rect 187262 18098 220706 18334
rect 220942 18098 221026 18334
rect 221262 18098 254706 18334
rect 254942 18098 255026 18334
rect 255262 18098 288706 18334
rect 288942 18098 289026 18334
rect 289262 18098 322706 18334
rect 322942 18098 323026 18334
rect 323262 18098 356706 18334
rect 356942 18098 357026 18334
rect 357262 18098 390706 18334
rect 390942 18098 391026 18334
rect 391262 18098 424706 18334
rect 424942 18098 425026 18334
rect 425262 18098 458706 18334
rect 458942 18098 459026 18334
rect 459262 18098 492706 18334
rect 492942 18098 493026 18334
rect 493262 18098 526706 18334
rect 526942 18098 527026 18334
rect 527262 18098 560706 18334
rect 560942 18098 561026 18334
rect 561262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 50706 18014
rect 50942 17778 51026 18014
rect 51262 17778 84706 18014
rect 84942 17778 85026 18014
rect 85262 17778 118706 18014
rect 118942 17778 119026 18014
rect 119262 17778 152706 18014
rect 152942 17778 153026 18014
rect 153262 17778 186706 18014
rect 186942 17778 187026 18014
rect 187262 17778 220706 18014
rect 220942 17778 221026 18014
rect 221262 17778 254706 18014
rect 254942 17778 255026 18014
rect 255262 17778 288706 18014
rect 288942 17778 289026 18014
rect 289262 17778 322706 18014
rect 322942 17778 323026 18014
rect 323262 17778 356706 18014
rect 356942 17778 357026 18014
rect 357262 17778 390706 18014
rect 390942 17778 391026 18014
rect 391262 17778 424706 18014
rect 424942 17778 425026 18014
rect 425262 17778 458706 18014
rect 458942 17778 459026 18014
rect 459262 17778 492706 18014
rect 492942 17778 493026 18014
rect 493262 17778 526706 18014
rect 526942 17778 527026 18014
rect 527262 17778 560706 18014
rect 560942 17778 561026 18014
rect 561262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 46986 14614
rect 47222 14378 47306 14614
rect 47542 14378 80986 14614
rect 81222 14378 81306 14614
rect 81542 14378 114986 14614
rect 115222 14378 115306 14614
rect 115542 14378 148986 14614
rect 149222 14378 149306 14614
rect 149542 14378 182986 14614
rect 183222 14378 183306 14614
rect 183542 14378 216986 14614
rect 217222 14378 217306 14614
rect 217542 14378 250986 14614
rect 251222 14378 251306 14614
rect 251542 14378 284986 14614
rect 285222 14378 285306 14614
rect 285542 14378 318986 14614
rect 319222 14378 319306 14614
rect 319542 14378 352986 14614
rect 353222 14378 353306 14614
rect 353542 14378 386986 14614
rect 387222 14378 387306 14614
rect 387542 14378 420986 14614
rect 421222 14378 421306 14614
rect 421542 14378 454986 14614
rect 455222 14378 455306 14614
rect 455542 14378 488986 14614
rect 489222 14378 489306 14614
rect 489542 14378 522986 14614
rect 523222 14378 523306 14614
rect 523542 14378 556986 14614
rect 557222 14378 557306 14614
rect 557542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 46986 14294
rect 47222 14058 47306 14294
rect 47542 14058 80986 14294
rect 81222 14058 81306 14294
rect 81542 14058 114986 14294
rect 115222 14058 115306 14294
rect 115542 14058 148986 14294
rect 149222 14058 149306 14294
rect 149542 14058 182986 14294
rect 183222 14058 183306 14294
rect 183542 14058 216986 14294
rect 217222 14058 217306 14294
rect 217542 14058 250986 14294
rect 251222 14058 251306 14294
rect 251542 14058 284986 14294
rect 285222 14058 285306 14294
rect 285542 14058 318986 14294
rect 319222 14058 319306 14294
rect 319542 14058 352986 14294
rect 353222 14058 353306 14294
rect 353542 14058 386986 14294
rect 387222 14058 387306 14294
rect 387542 14058 420986 14294
rect 421222 14058 421306 14294
rect 421542 14058 454986 14294
rect 455222 14058 455306 14294
rect 455542 14058 488986 14294
rect 489222 14058 489306 14294
rect 489542 14058 522986 14294
rect 523222 14058 523306 14294
rect 523542 14058 556986 14294
rect 557222 14058 557306 14294
rect 557542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 43266 10894
rect 43502 10658 43586 10894
rect 43822 10658 77266 10894
rect 77502 10658 77586 10894
rect 77822 10658 111266 10894
rect 111502 10658 111586 10894
rect 111822 10658 145266 10894
rect 145502 10658 145586 10894
rect 145822 10658 179266 10894
rect 179502 10658 179586 10894
rect 179822 10658 213266 10894
rect 213502 10658 213586 10894
rect 213822 10658 247266 10894
rect 247502 10658 247586 10894
rect 247822 10658 281266 10894
rect 281502 10658 281586 10894
rect 281822 10658 315266 10894
rect 315502 10658 315586 10894
rect 315822 10658 349266 10894
rect 349502 10658 349586 10894
rect 349822 10658 383266 10894
rect 383502 10658 383586 10894
rect 383822 10658 417266 10894
rect 417502 10658 417586 10894
rect 417822 10658 451266 10894
rect 451502 10658 451586 10894
rect 451822 10658 485266 10894
rect 485502 10658 485586 10894
rect 485822 10658 519266 10894
rect 519502 10658 519586 10894
rect 519822 10658 553266 10894
rect 553502 10658 553586 10894
rect 553822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 43266 10574
rect 43502 10338 43586 10574
rect 43822 10338 77266 10574
rect 77502 10338 77586 10574
rect 77822 10338 111266 10574
rect 111502 10338 111586 10574
rect 111822 10338 145266 10574
rect 145502 10338 145586 10574
rect 145822 10338 179266 10574
rect 179502 10338 179586 10574
rect 179822 10338 213266 10574
rect 213502 10338 213586 10574
rect 213822 10338 247266 10574
rect 247502 10338 247586 10574
rect 247822 10338 281266 10574
rect 281502 10338 281586 10574
rect 281822 10338 315266 10574
rect 315502 10338 315586 10574
rect 315822 10338 349266 10574
rect 349502 10338 349586 10574
rect 349822 10338 383266 10574
rect 383502 10338 383586 10574
rect 383822 10338 417266 10574
rect 417502 10338 417586 10574
rect 417822 10338 451266 10574
rect 451502 10338 451586 10574
rect 451822 10338 485266 10574
rect 485502 10338 485586 10574
rect 485822 10338 519266 10574
rect 519502 10338 519586 10574
rect 519822 10338 553266 10574
rect 553502 10338 553586 10574
rect 553822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 39546 7174
rect 39782 6938 39866 7174
rect 40102 6938 73546 7174
rect 73782 6938 73866 7174
rect 74102 6938 107546 7174
rect 107782 6938 107866 7174
rect 108102 6938 141546 7174
rect 141782 6938 141866 7174
rect 142102 6938 175546 7174
rect 175782 6938 175866 7174
rect 176102 6938 209546 7174
rect 209782 6938 209866 7174
rect 210102 6938 243546 7174
rect 243782 6938 243866 7174
rect 244102 6938 277546 7174
rect 277782 6938 277866 7174
rect 278102 6938 311546 7174
rect 311782 6938 311866 7174
rect 312102 6938 345546 7174
rect 345782 6938 345866 7174
rect 346102 6938 379546 7174
rect 379782 6938 379866 7174
rect 380102 6938 413546 7174
rect 413782 6938 413866 7174
rect 414102 6938 447546 7174
rect 447782 6938 447866 7174
rect 448102 6938 481546 7174
rect 481782 6938 481866 7174
rect 482102 6938 515546 7174
rect 515782 6938 515866 7174
rect 516102 6938 549546 7174
rect 549782 6938 549866 7174
rect 550102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 39546 6854
rect 39782 6618 39866 6854
rect 40102 6618 73546 6854
rect 73782 6618 73866 6854
rect 74102 6618 107546 6854
rect 107782 6618 107866 6854
rect 108102 6618 141546 6854
rect 141782 6618 141866 6854
rect 142102 6618 175546 6854
rect 175782 6618 175866 6854
rect 176102 6618 209546 6854
rect 209782 6618 209866 6854
rect 210102 6618 243546 6854
rect 243782 6618 243866 6854
rect 244102 6618 277546 6854
rect 277782 6618 277866 6854
rect 278102 6618 311546 6854
rect 311782 6618 311866 6854
rect 312102 6618 345546 6854
rect 345782 6618 345866 6854
rect 346102 6618 379546 6854
rect 379782 6618 379866 6854
rect 380102 6618 413546 6854
rect 413782 6618 413866 6854
rect 414102 6618 447546 6854
rect 447782 6618 447866 6854
rect 448102 6618 481546 6854
rect 481782 6618 481866 6854
rect 482102 6618 515546 6854
rect 515782 6618 515866 6854
rect 516102 6618 549546 6854
rect 549782 6618 549866 6854
rect 550102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 35826 3454
rect 36062 3218 36146 3454
rect 36382 3218 69826 3454
rect 70062 3218 70146 3454
rect 70382 3218 103826 3454
rect 104062 3218 104146 3454
rect 104382 3218 137826 3454
rect 138062 3218 138146 3454
rect 138382 3218 171826 3454
rect 172062 3218 172146 3454
rect 172382 3218 205826 3454
rect 206062 3218 206146 3454
rect 206382 3218 239826 3454
rect 240062 3218 240146 3454
rect 240382 3218 273826 3454
rect 274062 3218 274146 3454
rect 274382 3218 307826 3454
rect 308062 3218 308146 3454
rect 308382 3218 341826 3454
rect 342062 3218 342146 3454
rect 342382 3218 375826 3454
rect 376062 3218 376146 3454
rect 376382 3218 409826 3454
rect 410062 3218 410146 3454
rect 410382 3218 443826 3454
rect 444062 3218 444146 3454
rect 444382 3218 477826 3454
rect 478062 3218 478146 3454
rect 478382 3218 511826 3454
rect 512062 3218 512146 3454
rect 512382 3218 545826 3454
rect 546062 3218 546146 3454
rect 546382 3218 579826 3454
rect 580062 3218 580146 3454
rect 580382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 35826 3134
rect 36062 2898 36146 3134
rect 36382 2898 69826 3134
rect 70062 2898 70146 3134
rect 70382 2898 103826 3134
rect 104062 2898 104146 3134
rect 104382 2898 137826 3134
rect 138062 2898 138146 3134
rect 138382 2898 171826 3134
rect 172062 2898 172146 3134
rect 172382 2898 205826 3134
rect 206062 2898 206146 3134
rect 206382 2898 239826 3134
rect 240062 2898 240146 3134
rect 240382 2898 273826 3134
rect 274062 2898 274146 3134
rect 274382 2898 307826 3134
rect 308062 2898 308146 3134
rect 308382 2898 341826 3134
rect 342062 2898 342146 3134
rect 342382 2898 375826 3134
rect 376062 2898 376146 3134
rect 376382 2898 409826 3134
rect 410062 2898 410146 3134
rect 410382 2898 443826 3134
rect 444062 2898 444146 3134
rect 444382 2898 477826 3134
rect 478062 2898 478146 3134
rect 478382 2898 511826 3134
rect 512062 2898 512146 3134
rect 512382 2898 545826 3134
rect 546062 2898 546146 3134
rect 546382 2898 579826 3134
rect 580062 2898 580146 3134
rect 580382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 35826 -346
rect 36062 -582 36146 -346
rect 36382 -582 69826 -346
rect 70062 -582 70146 -346
rect 70382 -582 103826 -346
rect 104062 -582 104146 -346
rect 104382 -582 137826 -346
rect 138062 -582 138146 -346
rect 138382 -582 171826 -346
rect 172062 -582 172146 -346
rect 172382 -582 205826 -346
rect 206062 -582 206146 -346
rect 206382 -582 239826 -346
rect 240062 -582 240146 -346
rect 240382 -582 273826 -346
rect 274062 -582 274146 -346
rect 274382 -582 307826 -346
rect 308062 -582 308146 -346
rect 308382 -582 341826 -346
rect 342062 -582 342146 -346
rect 342382 -582 375826 -346
rect 376062 -582 376146 -346
rect 376382 -582 409826 -346
rect 410062 -582 410146 -346
rect 410382 -582 443826 -346
rect 444062 -582 444146 -346
rect 444382 -582 477826 -346
rect 478062 -582 478146 -346
rect 478382 -582 511826 -346
rect 512062 -582 512146 -346
rect 512382 -582 545826 -346
rect 546062 -582 546146 -346
rect 546382 -582 579826 -346
rect 580062 -582 580146 -346
rect 580382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 35826 -666
rect 36062 -902 36146 -666
rect 36382 -902 69826 -666
rect 70062 -902 70146 -666
rect 70382 -902 103826 -666
rect 104062 -902 104146 -666
rect 104382 -902 137826 -666
rect 138062 -902 138146 -666
rect 138382 -902 171826 -666
rect 172062 -902 172146 -666
rect 172382 -902 205826 -666
rect 206062 -902 206146 -666
rect 206382 -902 239826 -666
rect 240062 -902 240146 -666
rect 240382 -902 273826 -666
rect 274062 -902 274146 -666
rect 274382 -902 307826 -666
rect 308062 -902 308146 -666
rect 308382 -902 341826 -666
rect 342062 -902 342146 -666
rect 342382 -902 375826 -666
rect 376062 -902 376146 -666
rect 376382 -902 409826 -666
rect 410062 -902 410146 -666
rect 410382 -902 443826 -666
rect 444062 -902 444146 -666
rect 444382 -902 477826 -666
rect 478062 -902 478146 -666
rect 478382 -902 511826 -666
rect 512062 -902 512146 -666
rect 512382 -902 545826 -666
rect 546062 -902 546146 -666
rect 546382 -902 579826 -666
rect 580062 -902 580146 -666
rect 580382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 39546 -1306
rect 39782 -1542 39866 -1306
rect 40102 -1542 73546 -1306
rect 73782 -1542 73866 -1306
rect 74102 -1542 107546 -1306
rect 107782 -1542 107866 -1306
rect 108102 -1542 141546 -1306
rect 141782 -1542 141866 -1306
rect 142102 -1542 175546 -1306
rect 175782 -1542 175866 -1306
rect 176102 -1542 209546 -1306
rect 209782 -1542 209866 -1306
rect 210102 -1542 243546 -1306
rect 243782 -1542 243866 -1306
rect 244102 -1542 277546 -1306
rect 277782 -1542 277866 -1306
rect 278102 -1542 311546 -1306
rect 311782 -1542 311866 -1306
rect 312102 -1542 345546 -1306
rect 345782 -1542 345866 -1306
rect 346102 -1542 379546 -1306
rect 379782 -1542 379866 -1306
rect 380102 -1542 413546 -1306
rect 413782 -1542 413866 -1306
rect 414102 -1542 447546 -1306
rect 447782 -1542 447866 -1306
rect 448102 -1542 481546 -1306
rect 481782 -1542 481866 -1306
rect 482102 -1542 515546 -1306
rect 515782 -1542 515866 -1306
rect 516102 -1542 549546 -1306
rect 549782 -1542 549866 -1306
rect 550102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 39546 -1626
rect 39782 -1862 39866 -1626
rect 40102 -1862 73546 -1626
rect 73782 -1862 73866 -1626
rect 74102 -1862 107546 -1626
rect 107782 -1862 107866 -1626
rect 108102 -1862 141546 -1626
rect 141782 -1862 141866 -1626
rect 142102 -1862 175546 -1626
rect 175782 -1862 175866 -1626
rect 176102 -1862 209546 -1626
rect 209782 -1862 209866 -1626
rect 210102 -1862 243546 -1626
rect 243782 -1862 243866 -1626
rect 244102 -1862 277546 -1626
rect 277782 -1862 277866 -1626
rect 278102 -1862 311546 -1626
rect 311782 -1862 311866 -1626
rect 312102 -1862 345546 -1626
rect 345782 -1862 345866 -1626
rect 346102 -1862 379546 -1626
rect 379782 -1862 379866 -1626
rect 380102 -1862 413546 -1626
rect 413782 -1862 413866 -1626
rect 414102 -1862 447546 -1626
rect 447782 -1862 447866 -1626
rect 448102 -1862 481546 -1626
rect 481782 -1862 481866 -1626
rect 482102 -1862 515546 -1626
rect 515782 -1862 515866 -1626
rect 516102 -1862 549546 -1626
rect 549782 -1862 549866 -1626
rect 550102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 43266 -2266
rect 43502 -2502 43586 -2266
rect 43822 -2502 77266 -2266
rect 77502 -2502 77586 -2266
rect 77822 -2502 111266 -2266
rect 111502 -2502 111586 -2266
rect 111822 -2502 145266 -2266
rect 145502 -2502 145586 -2266
rect 145822 -2502 179266 -2266
rect 179502 -2502 179586 -2266
rect 179822 -2502 213266 -2266
rect 213502 -2502 213586 -2266
rect 213822 -2502 247266 -2266
rect 247502 -2502 247586 -2266
rect 247822 -2502 281266 -2266
rect 281502 -2502 281586 -2266
rect 281822 -2502 315266 -2266
rect 315502 -2502 315586 -2266
rect 315822 -2502 349266 -2266
rect 349502 -2502 349586 -2266
rect 349822 -2502 383266 -2266
rect 383502 -2502 383586 -2266
rect 383822 -2502 417266 -2266
rect 417502 -2502 417586 -2266
rect 417822 -2502 451266 -2266
rect 451502 -2502 451586 -2266
rect 451822 -2502 485266 -2266
rect 485502 -2502 485586 -2266
rect 485822 -2502 519266 -2266
rect 519502 -2502 519586 -2266
rect 519822 -2502 553266 -2266
rect 553502 -2502 553586 -2266
rect 553822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 43266 -2586
rect 43502 -2822 43586 -2586
rect 43822 -2822 77266 -2586
rect 77502 -2822 77586 -2586
rect 77822 -2822 111266 -2586
rect 111502 -2822 111586 -2586
rect 111822 -2822 145266 -2586
rect 145502 -2822 145586 -2586
rect 145822 -2822 179266 -2586
rect 179502 -2822 179586 -2586
rect 179822 -2822 213266 -2586
rect 213502 -2822 213586 -2586
rect 213822 -2822 247266 -2586
rect 247502 -2822 247586 -2586
rect 247822 -2822 281266 -2586
rect 281502 -2822 281586 -2586
rect 281822 -2822 315266 -2586
rect 315502 -2822 315586 -2586
rect 315822 -2822 349266 -2586
rect 349502 -2822 349586 -2586
rect 349822 -2822 383266 -2586
rect 383502 -2822 383586 -2586
rect 383822 -2822 417266 -2586
rect 417502 -2822 417586 -2586
rect 417822 -2822 451266 -2586
rect 451502 -2822 451586 -2586
rect 451822 -2822 485266 -2586
rect 485502 -2822 485586 -2586
rect 485822 -2822 519266 -2586
rect 519502 -2822 519586 -2586
rect 519822 -2822 553266 -2586
rect 553502 -2822 553586 -2586
rect 553822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 46986 -3226
rect 47222 -3462 47306 -3226
rect 47542 -3462 80986 -3226
rect 81222 -3462 81306 -3226
rect 81542 -3462 114986 -3226
rect 115222 -3462 115306 -3226
rect 115542 -3462 148986 -3226
rect 149222 -3462 149306 -3226
rect 149542 -3462 182986 -3226
rect 183222 -3462 183306 -3226
rect 183542 -3462 216986 -3226
rect 217222 -3462 217306 -3226
rect 217542 -3462 250986 -3226
rect 251222 -3462 251306 -3226
rect 251542 -3462 284986 -3226
rect 285222 -3462 285306 -3226
rect 285542 -3462 318986 -3226
rect 319222 -3462 319306 -3226
rect 319542 -3462 352986 -3226
rect 353222 -3462 353306 -3226
rect 353542 -3462 386986 -3226
rect 387222 -3462 387306 -3226
rect 387542 -3462 420986 -3226
rect 421222 -3462 421306 -3226
rect 421542 -3462 454986 -3226
rect 455222 -3462 455306 -3226
rect 455542 -3462 488986 -3226
rect 489222 -3462 489306 -3226
rect 489542 -3462 522986 -3226
rect 523222 -3462 523306 -3226
rect 523542 -3462 556986 -3226
rect 557222 -3462 557306 -3226
rect 557542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 46986 -3546
rect 47222 -3782 47306 -3546
rect 47542 -3782 80986 -3546
rect 81222 -3782 81306 -3546
rect 81542 -3782 114986 -3546
rect 115222 -3782 115306 -3546
rect 115542 -3782 148986 -3546
rect 149222 -3782 149306 -3546
rect 149542 -3782 182986 -3546
rect 183222 -3782 183306 -3546
rect 183542 -3782 216986 -3546
rect 217222 -3782 217306 -3546
rect 217542 -3782 250986 -3546
rect 251222 -3782 251306 -3546
rect 251542 -3782 284986 -3546
rect 285222 -3782 285306 -3546
rect 285542 -3782 318986 -3546
rect 319222 -3782 319306 -3546
rect 319542 -3782 352986 -3546
rect 353222 -3782 353306 -3546
rect 353542 -3782 386986 -3546
rect 387222 -3782 387306 -3546
rect 387542 -3782 420986 -3546
rect 421222 -3782 421306 -3546
rect 421542 -3782 454986 -3546
rect 455222 -3782 455306 -3546
rect 455542 -3782 488986 -3546
rect 489222 -3782 489306 -3546
rect 489542 -3782 522986 -3546
rect 523222 -3782 523306 -3546
rect 523542 -3782 556986 -3546
rect 557222 -3782 557306 -3546
rect 557542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 50706 -4186
rect 50942 -4422 51026 -4186
rect 51262 -4422 84706 -4186
rect 84942 -4422 85026 -4186
rect 85262 -4422 118706 -4186
rect 118942 -4422 119026 -4186
rect 119262 -4422 152706 -4186
rect 152942 -4422 153026 -4186
rect 153262 -4422 186706 -4186
rect 186942 -4422 187026 -4186
rect 187262 -4422 220706 -4186
rect 220942 -4422 221026 -4186
rect 221262 -4422 254706 -4186
rect 254942 -4422 255026 -4186
rect 255262 -4422 288706 -4186
rect 288942 -4422 289026 -4186
rect 289262 -4422 322706 -4186
rect 322942 -4422 323026 -4186
rect 323262 -4422 356706 -4186
rect 356942 -4422 357026 -4186
rect 357262 -4422 390706 -4186
rect 390942 -4422 391026 -4186
rect 391262 -4422 424706 -4186
rect 424942 -4422 425026 -4186
rect 425262 -4422 458706 -4186
rect 458942 -4422 459026 -4186
rect 459262 -4422 492706 -4186
rect 492942 -4422 493026 -4186
rect 493262 -4422 526706 -4186
rect 526942 -4422 527026 -4186
rect 527262 -4422 560706 -4186
rect 560942 -4422 561026 -4186
rect 561262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 50706 -4506
rect 50942 -4742 51026 -4506
rect 51262 -4742 84706 -4506
rect 84942 -4742 85026 -4506
rect 85262 -4742 118706 -4506
rect 118942 -4742 119026 -4506
rect 119262 -4742 152706 -4506
rect 152942 -4742 153026 -4506
rect 153262 -4742 186706 -4506
rect 186942 -4742 187026 -4506
rect 187262 -4742 220706 -4506
rect 220942 -4742 221026 -4506
rect 221262 -4742 254706 -4506
rect 254942 -4742 255026 -4506
rect 255262 -4742 288706 -4506
rect 288942 -4742 289026 -4506
rect 289262 -4742 322706 -4506
rect 322942 -4742 323026 -4506
rect 323262 -4742 356706 -4506
rect 356942 -4742 357026 -4506
rect 357262 -4742 390706 -4506
rect 390942 -4742 391026 -4506
rect 391262 -4742 424706 -4506
rect 424942 -4742 425026 -4506
rect 425262 -4742 458706 -4506
rect 458942 -4742 459026 -4506
rect 459262 -4742 492706 -4506
rect 492942 -4742 493026 -4506
rect 493262 -4742 526706 -4506
rect 526942 -4742 527026 -4506
rect 527262 -4742 560706 -4506
rect 560942 -4742 561026 -4506
rect 561262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 54426 -5146
rect 54662 -5382 54746 -5146
rect 54982 -5382 88426 -5146
rect 88662 -5382 88746 -5146
rect 88982 -5382 122426 -5146
rect 122662 -5382 122746 -5146
rect 122982 -5382 156426 -5146
rect 156662 -5382 156746 -5146
rect 156982 -5382 190426 -5146
rect 190662 -5382 190746 -5146
rect 190982 -5382 224426 -5146
rect 224662 -5382 224746 -5146
rect 224982 -5382 258426 -5146
rect 258662 -5382 258746 -5146
rect 258982 -5382 292426 -5146
rect 292662 -5382 292746 -5146
rect 292982 -5382 326426 -5146
rect 326662 -5382 326746 -5146
rect 326982 -5382 360426 -5146
rect 360662 -5382 360746 -5146
rect 360982 -5382 394426 -5146
rect 394662 -5382 394746 -5146
rect 394982 -5382 428426 -5146
rect 428662 -5382 428746 -5146
rect 428982 -5382 462426 -5146
rect 462662 -5382 462746 -5146
rect 462982 -5382 496426 -5146
rect 496662 -5382 496746 -5146
rect 496982 -5382 530426 -5146
rect 530662 -5382 530746 -5146
rect 530982 -5382 564426 -5146
rect 564662 -5382 564746 -5146
rect 564982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 54426 -5466
rect 54662 -5702 54746 -5466
rect 54982 -5702 88426 -5466
rect 88662 -5702 88746 -5466
rect 88982 -5702 122426 -5466
rect 122662 -5702 122746 -5466
rect 122982 -5702 156426 -5466
rect 156662 -5702 156746 -5466
rect 156982 -5702 190426 -5466
rect 190662 -5702 190746 -5466
rect 190982 -5702 224426 -5466
rect 224662 -5702 224746 -5466
rect 224982 -5702 258426 -5466
rect 258662 -5702 258746 -5466
rect 258982 -5702 292426 -5466
rect 292662 -5702 292746 -5466
rect 292982 -5702 326426 -5466
rect 326662 -5702 326746 -5466
rect 326982 -5702 360426 -5466
rect 360662 -5702 360746 -5466
rect 360982 -5702 394426 -5466
rect 394662 -5702 394746 -5466
rect 394982 -5702 428426 -5466
rect 428662 -5702 428746 -5466
rect 428982 -5702 462426 -5466
rect 462662 -5702 462746 -5466
rect 462982 -5702 496426 -5466
rect 496662 -5702 496746 -5466
rect 496982 -5702 530426 -5466
rect 530662 -5702 530746 -5466
rect 530982 -5702 564426 -5466
rect 564662 -5702 564746 -5466
rect 564982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 58146 -6106
rect 58382 -6342 58466 -6106
rect 58702 -6342 92146 -6106
rect 92382 -6342 92466 -6106
rect 92702 -6342 126146 -6106
rect 126382 -6342 126466 -6106
rect 126702 -6342 160146 -6106
rect 160382 -6342 160466 -6106
rect 160702 -6342 194146 -6106
rect 194382 -6342 194466 -6106
rect 194702 -6342 228146 -6106
rect 228382 -6342 228466 -6106
rect 228702 -6342 262146 -6106
rect 262382 -6342 262466 -6106
rect 262702 -6342 296146 -6106
rect 296382 -6342 296466 -6106
rect 296702 -6342 330146 -6106
rect 330382 -6342 330466 -6106
rect 330702 -6342 364146 -6106
rect 364382 -6342 364466 -6106
rect 364702 -6342 398146 -6106
rect 398382 -6342 398466 -6106
rect 398702 -6342 432146 -6106
rect 432382 -6342 432466 -6106
rect 432702 -6342 466146 -6106
rect 466382 -6342 466466 -6106
rect 466702 -6342 500146 -6106
rect 500382 -6342 500466 -6106
rect 500702 -6342 534146 -6106
rect 534382 -6342 534466 -6106
rect 534702 -6342 568146 -6106
rect 568382 -6342 568466 -6106
rect 568702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 58146 -6426
rect 58382 -6662 58466 -6426
rect 58702 -6662 92146 -6426
rect 92382 -6662 92466 -6426
rect 92702 -6662 126146 -6426
rect 126382 -6662 126466 -6426
rect 126702 -6662 160146 -6426
rect 160382 -6662 160466 -6426
rect 160702 -6662 194146 -6426
rect 194382 -6662 194466 -6426
rect 194702 -6662 228146 -6426
rect 228382 -6662 228466 -6426
rect 228702 -6662 262146 -6426
rect 262382 -6662 262466 -6426
rect 262702 -6662 296146 -6426
rect 296382 -6662 296466 -6426
rect 296702 -6662 330146 -6426
rect 330382 -6662 330466 -6426
rect 330702 -6662 364146 -6426
rect 364382 -6662 364466 -6426
rect 364702 -6662 398146 -6426
rect 398382 -6662 398466 -6426
rect 398702 -6662 432146 -6426
rect 432382 -6662 432466 -6426
rect 432702 -6662 466146 -6426
rect 466382 -6662 466466 -6426
rect 466702 -6662 500146 -6426
rect 500382 -6662 500466 -6426
rect 500702 -6662 534146 -6426
rect 534382 -6662 534466 -6426
rect 534702 -6662 568146 -6426
rect 568382 -6662 568466 -6426
rect 568702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 61866 -7066
rect 62102 -7302 62186 -7066
rect 62422 -7302 95866 -7066
rect 96102 -7302 96186 -7066
rect 96422 -7302 129866 -7066
rect 130102 -7302 130186 -7066
rect 130422 -7302 163866 -7066
rect 164102 -7302 164186 -7066
rect 164422 -7302 197866 -7066
rect 198102 -7302 198186 -7066
rect 198422 -7302 231866 -7066
rect 232102 -7302 232186 -7066
rect 232422 -7302 265866 -7066
rect 266102 -7302 266186 -7066
rect 266422 -7302 299866 -7066
rect 300102 -7302 300186 -7066
rect 300422 -7302 333866 -7066
rect 334102 -7302 334186 -7066
rect 334422 -7302 367866 -7066
rect 368102 -7302 368186 -7066
rect 368422 -7302 401866 -7066
rect 402102 -7302 402186 -7066
rect 402422 -7302 435866 -7066
rect 436102 -7302 436186 -7066
rect 436422 -7302 469866 -7066
rect 470102 -7302 470186 -7066
rect 470422 -7302 503866 -7066
rect 504102 -7302 504186 -7066
rect 504422 -7302 537866 -7066
rect 538102 -7302 538186 -7066
rect 538422 -7302 571866 -7066
rect 572102 -7302 572186 -7066
rect 572422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 61866 -7386
rect 62102 -7622 62186 -7386
rect 62422 -7622 95866 -7386
rect 96102 -7622 96186 -7386
rect 96422 -7622 129866 -7386
rect 130102 -7622 130186 -7386
rect 130422 -7622 163866 -7386
rect 164102 -7622 164186 -7386
rect 164422 -7622 197866 -7386
rect 198102 -7622 198186 -7386
rect 198422 -7622 231866 -7386
rect 232102 -7622 232186 -7386
rect 232422 -7622 265866 -7386
rect 266102 -7622 266186 -7386
rect 266422 -7622 299866 -7386
rect 300102 -7622 300186 -7386
rect 300422 -7622 333866 -7386
rect 334102 -7622 334186 -7386
rect 334422 -7622 367866 -7386
rect 368102 -7622 368186 -7386
rect 368422 -7622 401866 -7386
rect 402102 -7622 402186 -7386
rect 402422 -7622 435866 -7386
rect 436102 -7622 436186 -7386
rect 436422 -7622 469866 -7386
rect 470102 -7622 470186 -7386
rect 470422 -7622 503866 -7386
rect 504102 -7622 504186 -7386
rect 504422 -7622 537866 -7386
rect 538102 -7622 538186 -7386
rect 538422 -7622 571866 -7386
rect 572102 -7622 572186 -7386
rect 572422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 216400
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 116000 0 1 75000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 145914 0 1 174800
box -13000 -15200 17500 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 35794 -7654 36414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 69794 -7654 70414 223020 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 69794 232680 70414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 103794 -7654 104414 214340 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 103794 225660 104414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 137794 -7654 138414 74063 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 137794 163280 138414 185520 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 137794 225660 138414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 171794 -7654 172414 214340 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 171794 225660 172414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 205794 -7654 206414 214340 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 205794 225660 206414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 239794 -7654 240414 214340 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 239794 225660 240414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 273794 -7654 274414 214340 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 273794 225660 274414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 214340 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 307794 225660 308414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 341794 -7654 342414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 375794 -7654 376414 214340 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 375794 225660 376414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 409794 -7654 410414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 443794 -7654 444414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 477794 -7654 478414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 511794 -7654 512414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 545794 -7654 546414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 579794 -7654 580414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 36866 592650 37486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 70866 592650 71486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 104866 592650 105486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 138866 592650 139486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 172866 592650 173486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 206866 592650 207486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 240866 592650 241486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 274866 592650 275486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 342866 592650 343486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 376866 592650 377486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 410866 592650 411486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 444866 592650 445486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 478866 592650 479486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 512866 592650 513486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 546866 592650 547486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 580866 592650 581486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 648866 592650 649486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 682866 592650 683486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 43234 -7654 43854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 77234 -7654 77854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 77234 225660 77854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 111234 -7654 111854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 111234 225660 111854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 145234 -7654 145854 74063 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 145234 179075 145854 185520 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 145234 225660 145854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 179234 -7654 179854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 179234 225660 179854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 213234 -7654 213854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 213234 225660 213854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 247234 -7654 247854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 247234 225660 247854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 281234 -7654 281854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 315234 -7654 315854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 315234 225660 315854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 349234 -7654 349854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 349234 225660 349854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 383234 -7654 383854 214340 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 383234 225660 383854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 417234 -7654 417854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 451234 -7654 451854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 485234 -7654 485854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 519234 -7654 519854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 553234 -7654 553854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 44306 592650 44926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 78306 592650 78926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 112306 592650 112926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 146306 592650 146926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 180306 592650 180926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 214306 592650 214926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 248306 592650 248926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 282306 592650 282926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 316306 592650 316926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 350306 592650 350926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 384306 592650 384926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 418306 592650 418926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 452306 592650 452926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 486306 592650 486926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 520306 592650 520926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 554306 592650 554926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 588306 592650 588926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 656306 592650 656926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 690306 592650 690926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 50674 -7654 51294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 50674 225560 51294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 84674 -7654 85294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 84674 225660 85294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 118674 -7654 119294 74063 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 118674 134417 119294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 118674 225660 119294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 152674 -7654 153294 74063 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 152674 225660 153294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 186674 -7654 187294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 186674 225660 187294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 220674 -7654 221294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 254674 -7654 255294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 254674 225660 255294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 288674 -7654 289294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 288674 225660 289294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 322674 -7654 323294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 322674 225660 323294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 356674 -7654 357294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 356674 225660 357294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 390674 -7654 391294 214340 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 390674 225660 391294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 424674 -7654 425294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 458674 -7654 459294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 492674 -7654 493294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 526674 -7654 527294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 560674 -7654 561294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 51746 592650 52366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 85746 592650 86366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 119746 592650 120366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 153746 592650 154366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 187746 592650 188366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 221746 592650 222366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 255746 592650 256366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 289746 592650 290366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 323746 592650 324366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 357746 592650 358366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 391746 592650 392366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 425746 592650 426366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 459746 592650 460366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 493746 592650 494366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 527746 592650 528366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 561746 592650 562366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 595746 592650 596366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 663746 592650 664366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 697746 592650 698366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 58114 -7654 58734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 58114 225560 58734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 92114 -7654 92734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 92114 225660 92734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 126114 -7654 126734 74063 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 126114 134417 126734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 126114 225660 126734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 160114 -7654 160734 74063 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 160114 134417 160734 165832 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 160114 194880 160734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 194114 -7654 194734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 194114 225660 194734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 228114 -7654 228734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 228114 225660 228734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 262114 -7654 262734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 262114 225660 262734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 296114 -7654 296734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 296114 225660 296734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 330114 -7654 330734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 330114 225660 330734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 364114 -7654 364734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 364114 225660 364734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 398114 -7654 398734 214340 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 398114 225660 398734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 432114 -7654 432734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 466114 -7654 466734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 500114 -7654 500734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 534114 -7654 534734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 568114 -7654 568734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 59186 592650 59806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 93186 592650 93806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 127186 592650 127806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 161186 592650 161806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 195186 592650 195806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 229186 592650 229806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 263186 592650 263806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 297186 592650 297806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 331186 592650 331806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 365186 592650 365806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 399186 592650 399806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 433186 592650 433806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 467186 592650 467806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 501186 592650 501806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 535186 592650 535806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 569186 592650 569806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 603186 592650 603806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 671186 592650 671806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 54394 -7654 55014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 54394 225560 55014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 88394 -7654 89014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 88394 225660 89014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 122394 -7654 123014 74063 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 122394 134417 123014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 122394 225660 123014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 156394 -7654 157014 74063 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 156394 225660 157014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 190394 -7654 191014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 224394 -7654 225014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 224394 225660 225014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 258394 -7654 259014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 258394 225660 259014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 292394 -7654 293014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 292394 225660 293014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 326394 -7654 327014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 326394 225660 327014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 360394 -7654 361014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 360394 225660 361014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 394394 -7654 395014 214340 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 394394 225660 395014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 428394 -7654 429014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 462394 -7654 463014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 496394 -7654 497014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 530394 -7654 531014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564394 -7654 565014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 55466 592650 56086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 89466 592650 90086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 123466 592650 124086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 157466 592650 158086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 191466 592650 192086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 225466 592650 226086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 259466 592650 260086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 293466 592650 294086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 327466 592650 328086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 361466 592650 362086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 395466 592650 396086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 429466 592650 430086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 463466 592650 464086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 497466 592650 498086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 531466 592650 532086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565466 592650 566086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 599466 592650 600086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 667466 592650 668086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 61834 -7654 62454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 61834 225560 62454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 95834 -7654 96454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 95834 225660 96454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 129834 -7654 130454 74063 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 129834 134417 130454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 163834 -7654 164454 74063 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 163834 134417 164454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 163834 225660 164454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 197834 -7654 198454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 197834 225660 198454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 231834 -7654 232454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 231834 225660 232454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 265834 -7654 266454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 265834 225660 266454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 299834 -7654 300454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 299834 225660 300454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 333834 -7654 334454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 333834 225660 334454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 367834 -7654 368454 214340 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 367834 225660 368454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 401834 -7654 402454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 435834 -7654 436454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 469834 -7654 470454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 503834 -7654 504454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537834 -7654 538454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 571834 -7654 572454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 62906 592650 63526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 96906 592650 97526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 130906 592650 131526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 164906 592650 165526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 198906 592650 199526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 232906 592650 233526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 266906 592650 267526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 300906 592650 301526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 334906 592650 335526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 368906 592650 369526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 402906 592650 403526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 436906 592650 437526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 470906 592650 471526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 504906 592650 505526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538906 592650 539526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 572906 592650 573526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 606906 592650 607526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 674906 592650 675526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 39514 -7654 40134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 73514 -7654 74134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 73514 225660 74134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 107514 -7654 108134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 107514 225660 108134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 141514 -7654 142134 74063 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 141514 225660 142134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 175514 -7654 176134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 175514 225660 176134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 209514 -7654 210134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 209514 225660 210134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 243514 -7654 244134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 243514 225660 244134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 277514 -7654 278134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 277514 225660 278134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 311514 -7654 312134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 345514 -7654 346134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 345514 225660 346134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 379514 -7654 380134 214340 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 379514 225660 380134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 413514 -7654 414134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 447514 -7654 448134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 481514 -7654 482134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 515514 -7654 516134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 549514 -7654 550134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 40586 592650 41206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 74586 592650 75206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 108586 592650 109206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 142586 592650 143206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 176586 592650 177206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 210586 592650 211206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 244586 592650 245206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 278586 592650 279206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 312586 592650 313206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 346586 592650 347206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 380586 592650 381206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 414586 592650 415206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 448586 592650 449206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 482586 592650 483206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 516586 592650 517206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 550586 592650 551206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 584586 592650 585206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 652586 592650 653206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 686586 592650 687206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 46954 -7654 47574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 46954 225560 47574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 80954 -7654 81574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 80954 225660 81574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 114954 -7654 115574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 114954 225660 115574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 148954 -7654 149574 74063 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 148954 179075 149574 185520 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 148954 225660 149574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 182954 -7654 183574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 182954 225660 183574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 216954 -7654 217574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 216954 225660 217574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 250954 -7654 251574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 284954 -7654 285574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 284954 225660 285574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 318954 -7654 319574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 318954 225660 319574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 352954 -7654 353574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 352954 225660 353574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 386954 -7654 387574 214340 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 386954 225660 387574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 420954 -7654 421574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 454954 -7654 455574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 488954 -7654 489574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 522954 -7654 523574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 556954 -7654 557574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 48026 592650 48646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 82026 592650 82646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 116026 592650 116646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 150026 592650 150646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 184026 592650 184646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 218026 592650 218646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 252026 592650 252646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 286026 592650 286646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 320026 592650 320646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 354026 592650 354646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 388026 592650 388646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 422026 592650 422646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 456026 592650 456646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 490026 592650 490646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 524026 592650 524646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 558026 592650 558646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592026 592650 592646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 660026 592650 660646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 694026 592650 694646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 172264 105336 172264 105336 0 vccd1
rlabel via4 145704 180776 145704 180776 0 vccd2
rlabel via4 162334 188216 162334 188216 0 vdda1
rlabel via4 160584 161656 160584 161656 0 vdda2
rlabel via4 394864 225873 394864 225873 0 vssa1
rlabel metal5 291962 675216 291962 675216 0 vssa2
rlabel via4 175984 109056 175984 109056 0 vssd1
rlabel via4 149424 184496 149424 184496 0 vssd2
rlabel metal2 580198 444601 580198 444601 0 analog_io[3]
rlabel metal3 115023 133212 115023 133212 0 cmp
rlabel via3 139541 165172 139541 165172 0 cmp_out_c
rlabel metal2 178894 70380 178894 70380 0 io_in[0]
rlabel metal3 175812 92325 175812 92325 0 io_in[10]
rlabel metal3 175812 93753 175812 93753 0 io_in[11]
rlabel metal3 175812 95151 175812 95151 0 io_in[12]
rlabel metal3 175812 97085 175812 97085 0 io_in[13]
rlabel metal3 175812 98581 175812 98581 0 io_in[14]
rlabel metal3 175812 100077 175812 100077 0 io_in[15]
rlabel metal3 175812 101573 175812 101573 0 io_in[16]
rlabel metal3 175812 103069 175812 103069 0 io_in[17]
rlabel metal3 175812 104497 175812 104497 0 io_in[18]
rlabel metal3 347392 135116 347392 135116 0 io_in[19]
rlabel metal2 178802 62492 178802 62492 0 io_in[1]
rlabel metal3 59340 191692 59340 191692 0 io_in[20]
rlabel metal2 75302 289816 75302 289816 0 io_in[21]
rlabel metal2 45034 180438 45034 180438 0 io_in[22]
rlabel metal2 40526 422545 40526 422545 0 io_in[23]
rlabel metal3 175812 113103 175812 113103 0 io_in[24]
rlabel metal3 175812 114969 175812 114969 0 io_in[25]
rlabel metal3 175812 116465 175812 116465 0 io_in[26]
rlabel metal3 175812 117961 175812 117961 0 io_in[27]
rlabel metal3 175812 119457 175812 119457 0 io_in[28]
rlabel metal3 1970 423572 1970 423572 0 io_in[29]
rlabel metal3 175812 80561 175812 80561 0 io_in[2]
rlabel metal3 175812 122313 175812 122313 0 io_in[30]
rlabel metal3 175812 123877 175812 123877 0 io_in[31]
rlabel metal3 2016 267172 2016 267172 0 io_in[32]
rlabel metal3 1832 214948 1832 214948 0 io_in[33]
rlabel metal3 1832 162860 1832 162860 0 io_in[34]
rlabel metal3 175812 129657 175812 129657 0 io_in[35]
rlabel metal3 175812 131153 175812 131153 0 io_in[36]
rlabel metal3 175812 132551 175812 132551 0 io_in[37]
rlabel metal3 175812 82125 175812 82125 0 io_in[3]
rlabel metal3 175812 83621 175812 83621 0 io_in[4]
rlabel metal3 175812 85117 175812 85117 0 io_in[5]
rlabel metal3 175812 86545 175812 86545 0 io_in[6]
rlabel metal3 175812 87973 175812 87973 0 io_in[7]
rlabel metal3 175812 89469 175812 89469 0 io_in[8]
rlabel metal3 175812 90897 175812 90897 0 io_in[9]
rlabel metal3 581908 33116 581908 33116 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 580198 537319 580198 537319 0 io_oeb[11]
rlabel metal2 422970 331840 422970 331840 0 io_oeb[12]
rlabel metal3 581908 644028 581908 644028 0 io_oeb[13]
rlabel metal3 581954 697204 581954 697204 0 io_oeb[14]
rlabel metal2 527206 390058 527206 390058 0 io_oeb[15]
rlabel metal2 462346 389412 462346 389412 0 io_oeb[16]
rlabel metal2 397486 388902 397486 388902 0 io_oeb[17]
rlabel metal2 332534 701940 332534 701940 0 io_oeb[18]
rlabel metal1 153870 411298 153870 411298 0 io_oeb[19]
rlabel metal2 580198 72505 580198 72505 0 io_oeb[1]
rlabel metal1 115092 180710 115092 180710 0 io_oeb[20]
rlabel via1 56718 215917 56718 215917 0 io_oeb[21]
rlabel metal2 44850 148121 44850 148121 0 io_oeb[22]
rlabel metal3 118036 73032 118036 73032 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 1786 606084 1786 606084 0 io_oeb[25]
rlabel metal3 1832 553860 1832 553860 0 io_oeb[26]
rlabel metal3 1924 501772 1924 501772 0 io_oeb[27]
rlabel metal3 1556 449548 1556 449548 0 io_oeb[28]
rlabel metal3 1832 397460 1832 397460 0 io_oeb[29]
rlabel metal3 582000 112812 582000 112812 0 io_oeb[2]
rlabel metal3 1556 345372 1556 345372 0 io_oeb[30]
rlabel metal3 1832 293148 1832 293148 0 io_oeb[31]
rlabel metal3 1832 241060 1832 241060 0 io_oeb[32]
rlabel metal3 1740 188836 1740 188836 0 io_oeb[33]
rlabel metal3 1832 136748 1832 136748 0 io_oeb[34]
rlabel metal3 1832 84660 1832 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1556 6460 1556 6460 0 io_oeb[37]
rlabel metal3 582046 152660 582046 152660 0 io_oeb[3]
rlabel metal3 581954 192508 581954 192508 0 io_oeb[4]
rlabel metal3 582184 232356 582184 232356 0 io_oeb[5]
rlabel metal2 579646 272051 579646 272051 0 io_oeb[6]
rlabel metal2 579646 324785 579646 324785 0 io_oeb[7]
rlabel metal2 580198 378301 580198 378301 0 io_oeb[8]
rlabel metal2 580198 431103 580198 431103 0 io_oeb[9]
rlabel metal3 115345 75140 115345 75140 0 io_out[0]
rlabel metal3 114977 91052 114977 91052 0 io_out[10]
rlabel metal3 582092 524484 582092 524484 0 io_out[11]
rlabel metal3 582138 577660 582138 577660 0 io_out[12]
rlabel metal3 115928 95200 115928 95200 0 io_out[13]
rlabel metal3 115974 96696 115974 96696 0 io_out[14]
rlabel metal3 115851 98804 115851 98804 0 io_out[15]
rlabel metal3 116564 100009 116564 100009 0 io_out[16]
rlabel metal3 115805 101796 115805 101796 0 io_out[17]
rlabel metal3 115299 103156 115299 103156 0 io_out[18]
rlabel metal3 116196 104497 116196 104497 0 io_out[19]
rlabel metal3 115299 76636 115299 76636 0 io_out[1]
rlabel metal2 44942 403308 44942 403308 0 io_out[20]
rlabel metal2 45402 404056 45402 404056 0 io_out[21]
rlabel metal2 45126 167552 45126 167552 0 io_out[22]
rlabel metal2 24334 406973 24334 406973 0 io_out[23]
rlabel metal3 116196 111705 116196 111705 0 io_out[24]
rlabel metal3 116196 113103 116196 113103 0 io_out[25]
rlabel metal3 2016 566916 2016 566916 0 io_out[26]
rlabel metal3 116196 116669 116196 116669 0 io_out[27]
rlabel metal3 2660 462604 2660 462604 0 io_out[28]
rlabel metal3 116196 119593 116196 119593 0 io_out[29]
rlabel metal3 116564 78423 116564 78423 0 io_out[2]
rlabel metal3 116196 121021 116196 121021 0 io_out[30]
rlabel metal3 116196 122449 116196 122449 0 io_out[31]
rlabel metal2 22862 189108 22862 189108 0 io_out[32]
rlabel metal3 116196 125305 116196 125305 0 io_out[33]
rlabel metal3 1970 149804 1970 149804 0 io_out[34]
rlabel metal3 2062 97580 2062 97580 0 io_out[35]
rlabel metal3 2016 58548 2016 58548 0 io_out[36]
rlabel metal3 1970 19380 1970 19380 0 io_out[37]
rlabel metal3 115023 80852 115023 80852 0 io_out[3]
rlabel metal3 115253 82348 115253 82348 0 io_out[4]
rlabel metal3 115345 83708 115345 83708 0 io_out[5]
rlabel metal3 115207 85340 115207 85340 0 io_out[6]
rlabel metal3 115161 86836 115161 86836 0 io_out[7]
rlabel metal3 115115 88196 115115 88196 0 io_out[8]
rlabel metal3 115069 89692 115069 89692 0 io_out[9]
rlabel metal2 125902 1928 125902 1928 0 la_data_in[0]
rlabel metal2 480562 37067 480562 37067 0 la_data_in[100]
rlabel metal2 484058 37254 484058 37254 0 la_data_in[101]
rlabel metal2 487646 32970 487646 32970 0 la_data_in[102]
rlabel metal2 491142 32936 491142 32936 0 la_data_in[103]
rlabel metal3 326991 54468 326991 54468 0 la_data_in[104]
rlabel metal2 498226 2574 498226 2574 0 la_data_in[105]
rlabel metal2 501814 36455 501814 36455 0 la_data_in[106]
rlabel metal2 505402 36778 505402 36778 0 la_data_in[107]
rlabel metal2 508898 1928 508898 1928 0 la_data_in[108]
rlabel metal3 336789 55828 336789 55828 0 la_data_in[109]
rlabel metal2 161322 2115 161322 2115 0 la_data_in[10]
rlabel metal2 515982 37220 515982 37220 0 la_data_in[110]
rlabel metal2 519570 32256 519570 32256 0 la_data_in[111]
rlabel metal2 523066 31576 523066 31576 0 la_data_in[112]
rlabel metal2 526654 32919 526654 32919 0 la_data_in[113]
rlabel metal3 346265 57188 346265 57188 0 la_data_in[114]
rlabel metal2 533738 37186 533738 37186 0 la_data_in[115]
rlabel metal2 537234 37118 537234 37118 0 la_data_in[116]
rlabel metal2 540822 28788 540822 28788 0 la_data_in[117]
rlabel metal2 544410 29536 544410 29536 0 la_data_in[118]
rlabel metal3 355695 42092 355695 42092 0 la_data_in[119]
rlabel metal2 156722 20094 156722 20094 0 la_data_in[11]
rlabel metal2 551494 37152 551494 37152 0 la_data_in[120]
rlabel metal2 554990 37084 554990 37084 0 la_data_in[121]
rlabel metal2 558578 28108 558578 28108 0 la_data_in[122]
rlabel metal2 562074 25354 562074 25354 0 la_data_in[123]
rlabel metal2 565662 24623 565662 24623 0 la_data_in[124]
rlabel metal1 367862 53074 367862 53074 0 la_data_in[125]
rlabel metal1 369610 58650 369610 58650 0 la_data_in[126]
rlabel metal3 371381 47532 371381 47532 0 la_data_in[127]
rlabel metal2 168406 33072 168406 33072 0 la_data_in[12]
rlabel metal2 171994 31559 171994 31559 0 la_data_in[13]
rlabel metal2 175490 32239 175490 32239 0 la_data_in[14]
rlabel metal2 179078 37679 179078 37679 0 la_data_in[15]
rlabel metal2 178710 33694 178710 33694 0 la_data_in[16]
rlabel metal1 161184 53482 161184 53482 0 la_data_in[17]
rlabel metal2 189750 30879 189750 30879 0 la_data_in[18]
rlabel metal2 193246 28907 193246 28907 0 la_data_in[19]
rlabel metal2 129398 1928 129398 1928 0 la_data_in[1]
rlabel metal2 196834 37747 196834 37747 0 la_data_in[20]
rlabel metal2 200330 31712 200330 31712 0 la_data_in[21]
rlabel metal1 170660 50626 170660 50626 0 la_data_in[22]
rlabel metal1 172316 60214 172316 60214 0 la_data_in[23]
rlabel metal2 211002 28159 211002 28159 0 la_data_in[24]
rlabel metal2 214498 37611 214498 37611 0 la_data_in[25]
rlabel metal2 218086 37543 218086 37543 0 la_data_in[26]
rlabel metal2 221582 30930 221582 30930 0 la_data_in[27]
rlabel metal1 181930 57426 181930 57426 0 la_data_in[28]
rlabel metal2 228758 37815 228758 37815 0 la_data_in[29]
rlabel metal2 132986 21546 132986 21546 0 la_data_in[2]
rlabel metal2 232254 37271 232254 37271 0 la_data_in[30]
rlabel metal2 235842 37594 235842 37594 0 la_data_in[31]
rlabel metal1 189750 60146 189750 60146 0 la_data_in[32]
rlabel metal3 191521 54604 191521 54604 0 la_data_in[33]
rlabel metal3 193361 51884 193361 51884 0 la_data_in[34]
rlabel metal2 250010 37560 250010 37560 0 la_data_in[35]
rlabel metal2 253506 35962 253506 35962 0 la_data_in[36]
rlabel metal2 257094 2234 257094 2234 0 la_data_in[37]
rlabel metal2 260682 2200 260682 2200 0 la_data_in[38]
rlabel metal2 264178 2047 264178 2047 0 la_data_in[39]
rlabel metal2 136482 1894 136482 1894 0 la_data_in[3]
rlabel metal2 267766 37203 267766 37203 0 la_data_in[40]
rlabel metal2 271262 28856 271262 28856 0 la_data_in[41]
rlabel metal2 274850 27530 274850 27530 0 la_data_in[42]
rlabel metal3 210703 50388 210703 50388 0 la_data_in[43]
rlabel metal3 212589 49028 212589 49028 0 la_data_in[44]
rlabel metal2 285430 37526 285430 37526 0 la_data_in[45]
rlabel metal2 289018 35894 289018 35894 0 la_data_in[46]
rlabel metal2 292606 2132 292606 2132 0 la_data_in[47]
rlabel metal2 296102 1979 296102 1979 0 la_data_in[48]
rlabel metal2 299690 1911 299690 1911 0 la_data_in[49]
rlabel metal2 140070 8779 140070 8779 0 la_data_in[4]
rlabel metal2 303186 2166 303186 2166 0 la_data_in[50]
rlabel metal2 306774 36863 306774 36863 0 la_data_in[51]
rlabel metal2 310270 25456 310270 25456 0 la_data_in[52]
rlabel metal2 313858 28822 313858 28822 0 la_data_in[53]
rlabel metal3 231219 58684 231219 58684 0 la_data_in[54]
rlabel metal2 320942 37492 320942 37492 0 la_data_in[55]
rlabel metal1 235658 54638 235658 54638 0 la_data_in[56]
rlabel metal2 328026 26136 328026 26136 0 la_data_in[57]
rlabel metal2 331614 24011 331614 24011 0 la_data_in[58]
rlabel metal2 335110 23467 335110 23467 0 la_data_in[59]
rlabel metal2 143566 2574 143566 2574 0 la_data_in[5]
rlabel metal1 243524 60078 243524 60078 0 la_data_in[60]
rlabel metal1 245318 53346 245318 53346 0 la_data_in[61]
rlabel metal2 345782 24674 345782 24674 0 la_data_in[62]
rlabel metal2 349278 22583 349278 22583 0 la_data_in[63]
rlabel metal2 352866 21903 352866 21903 0 la_data_in[64]
rlabel metal2 356362 31644 356362 31644 0 la_data_in[65]
rlabel metal1 254794 55930 254794 55930 0 la_data_in[66]
rlabel metal1 256726 47702 256726 47702 0 la_data_in[67]
rlabel metal2 367034 25422 367034 25422 0 la_data_in[68]
rlabel metal2 370622 20543 370622 20543 0 la_data_in[69]
rlabel metal1 134780 52462 134780 52462 0 la_data_in[6]
rlabel metal2 374118 30896 374118 30896 0 la_data_in[70]
rlabel metal1 264454 51850 264454 51850 0 la_data_in[71]
rlabel metal1 266156 60010 266156 60010 0 la_data_in[72]
rlabel metal2 384790 23399 384790 23399 0 la_data_in[73]
rlabel metal2 388286 19795 388286 19795 0 la_data_in[74]
rlabel metal2 391874 35826 391874 35826 0 la_data_in[75]
rlabel metal2 395370 37135 395370 37135 0 la_data_in[76]
rlabel metal1 275862 44982 275862 44982 0 la_data_in[77]
rlabel metal1 277702 42126 277702 42126 0 la_data_in[78]
rlabel metal2 406042 19115 406042 19115 0 la_data_in[79]
rlabel metal2 150650 1962 150650 1962 0 la_data_in[7]
rlabel metal2 409630 29570 409630 29570 0 la_data_in[80]
rlabel metal1 283590 53278 283590 53278 0 la_data_in[81]
rlabel metal1 285430 47634 285430 47634 0 la_data_in[82]
rlabel metal3 287063 40596 287063 40596 0 la_data_in[83]
rlabel metal2 423798 18435 423798 18435 0 la_data_in[84]
rlabel metal2 427294 27462 427294 27462 0 la_data_in[85]
rlabel metal2 430882 25388 430882 25388 0 la_data_in[86]
rlabel metal1 294906 43554 294906 43554 0 la_data_in[87]
rlabel metal3 296677 51748 296677 51748 0 la_data_in[88]
rlabel metal3 298563 35292 298563 35292 0 la_data_in[89]
rlabel metal2 154238 1928 154238 1928 0 la_data_in[8]
rlabel metal2 445050 36472 445050 36472 0 la_data_in[90]
rlabel metal2 448638 35792 448638 35792 0 la_data_in[91]
rlabel metal2 452134 2064 452134 2064 0 la_data_in[92]
rlabel metal2 455722 1996 455722 1996 0 la_data_in[93]
rlabel metal2 459218 1843 459218 1843 0 la_data_in[94]
rlabel metal2 462806 2030 462806 2030 0 la_data_in[95]
rlabel metal2 466302 35078 466302 35078 0 la_data_in[96]
rlabel metal2 469890 35044 469890 35044 0 la_data_in[97]
rlabel metal2 473478 3339 473478 3339 0 la_data_in[98]
rlabel metal2 476974 3271 476974 3271 0 la_data_in[99]
rlabel metal2 157826 1928 157826 1928 0 la_data_in[9]
rlabel metal2 127006 1894 127006 1894 0 la_data_out[0]
rlabel metal2 481758 21920 481758 21920 0 la_data_out[100]
rlabel metal2 485254 15766 485254 15766 0 la_data_out[101]
rlabel metal2 488842 14338 488842 14338 0 la_data_out[102]
rlabel metal3 325887 26860 325887 26860 0 la_data_out[103]
rlabel metal1 328532 35190 328532 35190 0 la_data_out[104]
rlabel metal1 330188 40698 330188 40698 0 la_data_out[105]
rlabel metal2 503010 12978 503010 12978 0 la_data_out[106]
rlabel metal2 506506 19880 506506 19880 0 la_data_out[107]
rlabel metal1 335386 24174 335386 24174 0 la_data_out[108]
rlabel metal1 337548 22746 337548 22746 0 la_data_out[109]
rlabel metal2 160770 22338 160770 22338 0 la_data_out[10]
rlabel metal1 339802 33762 339802 33762 0 la_data_out[110]
rlabel metal2 520766 16378 520766 16378 0 la_data_out[111]
rlabel metal2 524262 1962 524262 1962 0 la_data_out[112]
rlabel metal2 527850 5991 527850 5991 0 la_data_out[113]
rlabel metal1 347714 8942 347714 8942 0 la_data_out[114]
rlabel metal1 349462 10302 349462 10302 0 la_data_out[115]
rlabel metal2 538430 35724 538430 35724 0 la_data_out[116]
rlabel metal2 542018 3968 542018 3968 0 la_data_out[117]
rlabel metal2 545514 35690 545514 35690 0 la_data_out[118]
rlabel metal1 357190 31042 357190 31042 0 la_data_out[119]
rlabel metal1 138115 3366 138115 3366 0 la_data_out[11]
rlabel metal1 358892 53142 358892 53142 0 la_data_out[120]
rlabel metal2 556186 3288 556186 3288 0 la_data_out[121]
rlabel metal2 559774 35707 559774 35707 0 la_data_out[122]
rlabel metal2 563270 14967 563270 14967 0 la_data_out[123]
rlabel metal2 566858 14304 566858 14304 0 la_data_out[124]
rlabel metal1 368138 26894 368138 26894 0 la_data_out[125]
rlabel metal1 370300 37910 370300 37910 0 la_data_out[126]
rlabel metal2 577438 6671 577438 6671 0 la_data_out[127]
rlabel metal2 169602 34840 169602 34840 0 la_data_out[12]
rlabel metal2 135010 74725 135010 74725 0 la_data_out[13]
rlabel metal2 176686 29638 176686 29638 0 la_data_out[14]
rlabel metal2 180274 24096 180274 24096 0 la_data_out[15]
rlabel metal1 159804 39542 159804 39542 0 la_data_out[16]
rlabel metal2 187358 2098 187358 2098 0 la_data_out[17]
rlabel metal2 190854 19863 190854 19863 0 la_data_out[18]
rlabel metal2 194442 35622 194442 35622 0 la_data_out[19]
rlabel metal2 130594 1894 130594 1894 0 la_data_out[1]
rlabel metal2 197938 21988 197938 21988 0 la_data_out[20]
rlabel metal1 169418 53414 169418 53414 0 la_data_out[21]
rlabel metal2 205114 3220 205114 3220 0 la_data_out[22]
rlabel metal2 208610 35775 208610 35775 0 la_data_out[23]
rlabel metal2 212198 21308 212198 21308 0 la_data_out[24]
rlabel metal2 215694 20628 215694 20628 0 la_data_out[25]
rlabel metal2 219282 16514 219282 16514 0 la_data_out[26]
rlabel metal1 180642 16150 180642 16150 0 la_data_out[27]
rlabel metal3 182781 25636 182781 25636 0 la_data_out[28]
rlabel metal2 229862 1860 229862 1860 0 la_data_out[29]
rlabel metal2 134037 340 134037 340 0 la_data_out[2]
rlabel metal2 233450 15834 233450 15834 0 la_data_out[30]
rlabel metal2 237038 12400 237038 12400 0 la_data_out[31]
rlabel metal1 190210 13362 190210 13362 0 la_data_out[32]
rlabel metal3 192303 36652 192303 36652 0 la_data_out[33]
rlabel metal2 247618 35656 247618 35656 0 la_data_out[34]
rlabel metal2 251206 35996 251206 35996 0 la_data_out[35]
rlabel metal2 254702 3526 254702 3526 0 la_data_out[36]
rlabel metal2 258290 3492 258290 3492 0 la_data_out[37]
rlabel metal2 261786 3458 261786 3458 0 la_data_out[38]
rlabel metal1 203780 7786 203780 7786 0 la_data_out[39]
rlabel metal2 137678 3288 137678 3288 0 la_data_out[3]
rlabel metal2 268870 14440 268870 14440 0 la_data_out[40]
rlabel metal2 272458 17874 272458 17874 0 la_data_out[41]
rlabel metal2 276046 7538 276046 7538 0 la_data_out[42]
rlabel metal2 279542 32307 279542 32307 0 la_data_out[43]
rlabel metal2 283130 35928 283130 35928 0 la_data_out[44]
rlabel metal1 215234 39474 215234 39474 0 la_data_out[45]
rlabel metal2 290214 7504 290214 7504 0 la_data_out[46]
rlabel metal2 293710 16480 293710 16480 0 la_data_out[47]
rlabel metal3 220823 9044 220823 9044 0 la_data_out[48]
rlabel metal1 223284 38046 223284 38046 0 la_data_out[49]
rlabel metal2 141266 1656 141266 1656 0 la_data_out[4]
rlabel metal1 225124 25738 225124 25738 0 la_data_out[50]
rlabel metal2 307970 35860 307970 35860 0 la_data_out[51]
rlabel metal2 311466 35282 311466 35282 0 la_data_out[52]
rlabel metal2 315054 13726 315054 13726 0 la_data_out[53]
rlabel metal1 232852 24378 232852 24378 0 la_data_out[54]
rlabel metal2 322138 2710 322138 2710 0 la_data_out[55]
rlabel metal1 236486 13294 236486 13294 0 la_data_out[56]
rlabel metal2 329222 5430 329222 5430 0 la_data_out[57]
rlabel metal2 332718 11567 332718 11567 0 la_data_out[58]
rlabel metal1 242236 14586 242236 14586 0 la_data_out[59]
rlabel metal1 139104 43418 139104 43418 0 la_data_out[5]
rlabel metal1 243938 7718 243938 7718 0 la_data_out[60]
rlabel metal2 343390 37458 343390 37458 0 la_data_out[61]
rlabel metal2 346978 2098 346978 2098 0 la_data_out[62]
rlabel metal2 350474 5311 350474 5311 0 la_data_out[63]
rlabel metal2 354062 35248 354062 35248 0 la_data_out[64]
rlabel metal1 253828 31246 253828 31246 0 la_data_out[65]
rlabel metal1 255576 42194 255576 42194 0 la_data_out[66]
rlabel metal2 364642 4750 364642 4750 0 la_data_out[67]
rlabel metal2 368230 34959 368230 34959 0 la_data_out[68]
rlabel metal2 371726 13012 371726 13012 0 la_data_out[69]
rlabel metal1 140990 21386 140990 21386 0 la_data_out[6]
rlabel metal1 263028 16014 263028 16014 0 la_data_out[70]
rlabel metal1 264730 15946 264730 15946 0 la_data_out[71]
rlabel metal2 382398 35214 382398 35214 0 la_data_out[72]
rlabel metal2 385986 6059 385986 6059 0 la_data_out[73]
rlabel metal2 389482 12332 389482 12332 0 la_data_out[74]
rlabel metal2 393070 8116 393070 8116 0 la_data_out[75]
rlabel metal2 396566 35180 396566 35180 0 la_data_out[76]
rlabel metal2 400154 2608 400154 2608 0 la_data_out[77]
rlabel metal2 403650 35146 403650 35146 0 la_data_out[78]
rlabel metal2 407238 35112 407238 35112 0 la_data_out[79]
rlabel metal2 151846 3254 151846 3254 0 la_data_out[7]
rlabel metal2 410826 6790 410826 6790 0 la_data_out[80]
rlabel metal1 284280 14450 284280 14450 0 la_data_out[81]
rlabel metal2 417910 3356 417910 3356 0 la_data_out[82]
rlabel metal3 287845 22644 287845 22644 0 la_data_out[83]
rlabel metal2 424994 17092 424994 17092 0 la_data_out[84]
rlabel metal2 428490 4002 428490 4002 0 la_data_out[85]
rlabel metal1 293756 36550 293756 36550 0 la_data_out[86]
rlabel metal1 295642 10438 295642 10438 0 la_data_out[87]
rlabel metal3 297183 59908 297183 59908 0 la_data_out[88]
rlabel metal2 442658 23960 442658 23960 0 la_data_out[89]
rlabel metal2 155434 1996 155434 1996 0 la_data_out[8]
rlabel metal2 446246 33004 446246 33004 0 la_data_out[90]
rlabel metal2 449834 14372 449834 14372 0 la_data_out[91]
rlabel metal2 453330 30862 453330 30862 0 la_data_out[92]
rlabel metal3 306521 35156 306521 35156 0 la_data_out[93]
rlabel metal1 308890 29614 308890 29614 0 la_data_out[94]
rlabel metal2 464002 8864 464002 8864 0 la_data_out[95]
rlabel metal2 467498 8830 467498 8830 0 la_data_out[96]
rlabel metal1 314456 17238 314456 17238 0 la_data_out[97]
rlabel metal3 316181 57324 316181 57324 0 la_data_out[98]
rlabel metal1 318688 9010 318688 9010 0 la_data_out[99]
rlabel metal2 158930 1826 158930 1826 0 la_data_out[9]
rlabel metal2 131514 73450 131514 73450 0 la_oenb[0]
rlabel metal2 482862 6042 482862 6042 0 la_oenb[100]
rlabel metal2 486450 20560 486450 20560 0 la_oenb[101]
rlabel metal3 324783 15844 324783 15844 0 la_oenb[102]
rlabel metal2 493534 2591 493534 2591 0 la_oenb[103]
rlabel metal2 497122 35010 497122 35010 0 la_oenb[104]
rlabel metal2 500618 22600 500618 22600 0 la_oenb[105]
rlabel metal2 504206 35758 504206 35758 0 la_oenb[106]
rlabel metal2 507702 13658 507702 13658 0 la_oenb[107]
rlabel metal3 336283 50252 336283 50252 0 la_oenb[108]
rlabel metal1 338514 43418 338514 43418 0 la_oenb[109]
rlabel metal2 163714 1928 163714 1928 0 la_oenb[10]
rlabel metal1 340492 32470 340492 32470 0 la_oenb[110]
rlabel metal2 521870 12944 521870 12944 0 la_oenb[111]
rlabel metal2 525458 21206 525458 21206 0 la_oenb[112]
rlabel metal3 345805 14484 345805 14484 0 la_oenb[113]
rlabel metal1 348220 24106 348220 24106 0 la_oenb[114]
rlabel metal1 349968 31110 349968 31110 0 la_oenb[115]
rlabel metal2 539626 26782 539626 26782 0 la_oenb[116]
rlabel metal2 543214 19846 543214 19846 0 la_oenb[117]
rlabel metal2 546710 1996 546710 1996 0 la_oenb[118]
rlabel metal1 357834 13090 357834 13090 0 la_oenb[119]
rlabel metal2 167210 34602 167210 34602 0 la_oenb[11]
rlabel metal2 553794 34432 553794 34432 0 la_oenb[120]
rlabel metal2 557382 3254 557382 3254 0 la_oenb[121]
rlabel metal2 560878 34398 560878 34398 0 la_oenb[122]
rlabel metal2 564466 9527 564466 9527 0 la_oenb[123]
rlabel metal2 568054 34364 568054 34364 0 la_oenb[124]
rlabel metal1 368828 18598 368828 18598 0 la_oenb[125]
rlabel metal2 575138 34330 575138 34330 0 la_oenb[126]
rlabel metal2 578634 9459 578634 9459 0 la_oenb[127]
rlabel metal2 170798 34483 170798 34483 0 la_oenb[12]
rlabel metal2 174294 26187 174294 26187 0 la_oenb[13]
rlabel metal2 177882 28176 177882 28176 0 la_oenb[14]
rlabel metal2 181470 34568 181470 34568 0 la_oenb[15]
rlabel metal1 160632 49062 160632 49062 0 la_oenb[16]
rlabel metal1 162104 46274 162104 46274 0 la_oenb[17]
rlabel metal2 192050 34415 192050 34415 0 la_oenb[18]
rlabel metal2 195638 3186 195638 3186 0 la_oenb[19]
rlabel metal1 131790 65212 131790 65212 0 la_oenb[1]
rlabel metal2 199134 2744 199134 2744 0 la_oenb[20]
rlabel metal1 170200 18802 170200 18802 0 la_oenb[21]
rlabel metal1 171902 38114 171902 38114 0 la_oenb[22]
rlabel metal2 209806 13675 209806 13675 0 la_oenb[23]
rlabel metal2 213394 34534 213394 34534 0 la_oenb[24]
rlabel metal2 216890 27564 216890 27564 0 la_oenb[25]
rlabel metal1 179400 17510 179400 17510 0 la_oenb[26]
rlabel metal1 181562 28594 181562 28594 0 la_oenb[27]
rlabel metal2 227562 34347 227562 34347 0 la_oenb[28]
rlabel metal2 231058 11006 231058 11006 0 la_oenb[29]
rlabel metal2 135286 1928 135286 1928 0 la_oenb[2]
rlabel metal2 234646 23280 234646 23280 0 la_oenb[30]
rlabel metal2 238142 9544 238142 9544 0 la_oenb[31]
rlabel metal2 241730 34500 241730 34500 0 la_oenb[32]
rlabel metal3 192947 11900 192947 11900 0 la_oenb[33]
rlabel metal2 248814 3594 248814 3594 0 la_oenb[34]
rlabel metal2 252402 3560 252402 3560 0 la_oenb[35]
rlabel metal2 255898 3407 255898 3407 0 la_oenb[36]
rlabel metal1 200468 36686 200468 36686 0 la_oenb[37]
rlabel metal2 262982 35027 262982 35027 0 la_oenb[38]
rlabel metal1 204930 20230 204930 20230 0 la_oenb[39]
rlabel metal2 138874 1843 138874 1843 0 la_oenb[3]
rlabel metal2 270066 20594 270066 20594 0 la_oenb[40]
rlabel metal2 273654 17126 273654 17126 0 la_oenb[41]
rlabel metal2 277150 29604 277150 29604 0 la_oenb[42]
rlabel metal3 211807 19924 211807 19924 0 la_oenb[43]
rlabel metal1 214452 20162 214452 20162 0 la_oenb[44]
rlabel metal2 287822 11618 287822 11618 0 la_oenb[45]
rlabel metal2 291410 24062 291410 24062 0 la_oenb[46]
rlabel metal2 294906 10224 294906 10224 0 la_oenb[47]
rlabel metal2 298494 33667 298494 33667 0 la_oenb[48]
rlabel metal2 301990 3424 301990 3424 0 la_oenb[49]
rlabel metal1 138000 32402 138000 32402 0 la_oenb[4]
rlabel metal2 305578 3390 305578 3390 0 la_oenb[50]
rlabel metal2 309074 4818 309074 4818 0 la_oenb[51]
rlabel metal2 312662 4784 312662 4784 0 la_oenb[52]
rlabel metal3 231219 8908 231219 8908 0 la_oenb[53]
rlabel metal1 233404 35326 233404 35326 0 la_oenb[54]
rlabel metal1 235290 16082 235290 16082 0 la_oenb[55]
rlabel metal2 326830 33718 326830 33718 0 la_oenb[56]
rlabel metal2 330418 2676 330418 2676 0 la_oenb[57]
rlabel metal2 333914 33599 333914 33599 0 la_oenb[58]
rlabel metal1 243064 32538 243064 32538 0 la_oenb[59]
rlabel metal2 145958 2030 145958 2030 0 la_oenb[5]
rlabel metal1 244904 21590 244904 21590 0 la_oenb[60]
rlabel metal1 246652 21522 246652 21522 0 la_oenb[61]
rlabel metal2 348082 33684 348082 33684 0 la_oenb[62]
rlabel metal2 351670 10819 351670 10819 0 la_oenb[63]
rlabel metal2 355258 33650 355258 33650 0 la_oenb[64]
rlabel metal1 253966 21454 253966 21454 0 la_oenb[65]
rlabel metal1 258106 37978 258106 37978 0 la_oenb[66]
rlabel metal2 365838 10870 365838 10870 0 la_oenb[67]
rlabel metal2 369426 33616 369426 33616 0 la_oenb[68]
rlabel metal2 372922 14406 372922 14406 0 la_oenb[69]
rlabel metal2 149546 1996 149546 1996 0 la_oenb[6]
rlabel metal1 264040 18666 264040 18666 0 la_oenb[70]
rlabel metal1 265696 27030 265696 27030 0 la_oenb[71]
rlabel metal1 271492 20026 271492 20026 0 la_oenb[72]
rlabel metal2 387182 17075 387182 17075 0 la_oenb[73]
rlabel metal2 390678 2642 390678 2642 0 la_oenb[74]
rlabel metal2 394266 31610 394266 31610 0 la_oenb[75]
rlabel metal2 397762 32290 397762 32290 0 la_oenb[76]
rlabel metal1 284740 22814 284740 22814 0 la_oenb[77]
rlabel metal2 404846 12927 404846 12927 0 la_oenb[78]
rlabel metal2 408434 12298 408434 12298 0 la_oenb[79]
rlabel metal2 153042 2166 153042 2166 0 la_oenb[7]
rlabel metal2 411930 4716 411930 4716 0 la_oenb[80]
rlabel metal1 291686 11798 291686 11798 0 la_oenb[81]
rlabel metal3 286741 7548 286741 7548 0 la_oenb[82]
rlabel metal2 422602 7436 422602 7436 0 la_oenb[83]
rlabel metal2 426190 6756 426190 6756 0 la_oenb[84]
rlabel metal2 429686 18486 429686 18486 0 la_oenb[85]
rlabel metal2 433274 3322 433274 3322 0 la_oenb[86]
rlabel metal1 302174 51782 302174 51782 0 la_oenb[87]
rlabel metal3 298057 30940 298057 30940 0 la_oenb[88]
rlabel metal2 443854 8898 443854 8898 0 la_oenb[89]
rlabel metal2 156630 21223 156630 21223 0 la_oenb[8]
rlabel metal2 447442 22634 447442 22634 0 la_oenb[90]
rlabel metal2 450938 10156 450938 10156 0 la_oenb[91]
rlabel metal1 305762 29682 305762 29682 0 la_oenb[92]
rlabel metal2 169050 37615 169050 37615 0 la_oenb[93]
rlabel metal2 461610 34466 461610 34466 0 la_oenb[94]
rlabel metal2 465198 17806 465198 17806 0 la_oenb[95]
rlabel metal2 468694 27428 468694 27428 0 la_oenb[96]
rlabel metal2 332626 69887 332626 69887 0 la_oenb[97]
rlabel metal2 173282 35343 173282 35343 0 la_oenb[98]
rlabel metal1 475318 8262 475318 8262 0 la_oenb[99]
rlabel metal2 160126 1656 160126 1656 0 la_oenb[9]
rlabel metal2 156906 136330 156906 136330 0 ota_out_c
rlabel metal3 151133 152388 151133 152388 0 ota_sh_c
rlabel metal2 57829 214540 57829 214540 0 pd1
rlabel metal2 327106 199369 327106 199369 0 pd10
rlabel metal3 135608 160004 135608 160004 0 pd10_a
rlabel metal2 124062 136466 124062 136466 0 pd10_b
rlabel metal3 355948 212636 355948 212636 0 pd11
rlabel metal2 122498 136211 122498 136211 0 pd11_a
rlabel metal2 121125 134980 121125 134980 0 pd11_b
rlabel metal2 386538 213853 386538 213853 0 pd12
rlabel metal2 119370 135990 119370 135990 0 pd12_a
rlabel metal2 117997 134980 117997 134980 0 pd12_b
rlabel metal2 153778 136432 153778 136432 0 pd1_a
rlabel metal2 152214 136398 152214 136398 0 pd1_b
rlabel via2 133262 182019 133262 182019 0 pd2
rlabel metal2 150650 135990 150650 135990 0 pd2_a
rlabel metal2 149086 135888 149086 135888 0 pd2_b
rlabel metal2 133262 180047 133262 180047 0 pd3
rlabel metal2 147522 136466 147522 136466 0 pd3_a
rlabel metal2 145767 134980 145767 134980 0 pd3_b
rlabel metal2 146411 214540 146411 214540 0 pd4
rlabel metal2 144295 134980 144295 134980 0 pd4_a
rlabel metal2 142830 147356 142830 147356 0 pd4_b
rlabel metal1 175628 211106 175628 211106 0 pd5
rlabel metal2 141365 134980 141365 134980 0 pd5_a
rlabel metal2 139893 134980 139893 134980 0 pd5_b
rlabel metal1 176640 188326 176640 188326 0 pd6
rlabel metal2 138375 134980 138375 134980 0 pd6_a
rlabel metal1 137632 157386 137632 157386 0 pd6_b
rlabel metal2 236295 214540 236295 214540 0 pd7
rlabel metal2 135010 136432 135010 136432 0 pd7_a
rlabel metal2 133637 134980 133637 134980 0 pd7_b
rlabel metal1 207966 191114 207966 191114 0 pd8
rlabel metal2 135654 158892 135654 158892 0 pd8_a
rlabel metal2 134550 158552 134550 158552 0 pd8_b
rlabel metal2 296746 213853 296746 213853 0 pd9
rlabel via2 136390 179469 136390 179469 0 pd9_a
rlabel metal2 127381 134980 127381 134980 0 pd9_b
rlabel metal2 174011 134980 174011 134980 0 sh
rlabel metal2 172546 136126 172546 136126 0 sh_cmp
rlabel metal2 158470 136058 158470 136058 0 sh_out_c
rlabel metal2 170982 136160 170982 136160 0 sh_rst
rlabel metal2 169227 134980 169227 134980 0 sw1
rlabel metal2 167854 136211 167854 136211 0 sw2
rlabel metal2 581026 23263 581026 23263 0 user_irq[0]
rlabel metal2 582222 1826 582222 1826 0 user_irq[1]
rlabel metal2 583418 1894 583418 1894 0 user_irq[2]
rlabel metal1 149546 161262 149546 161262 0 vd1
rlabel metal2 166099 134980 166099 134980 0 vd2
rlabel metal2 160034 135854 160034 135854 0 vref_cmp_c
rlabel metal2 155342 136466 155342 136466 0 vref_sel_c
rlabel metal2 598 1894 598 1894 0 wb_clk_i
rlabel metal2 1702 1928 1702 1928 0 wb_rst_i
rlabel metal2 2898 32936 2898 32936 0 wbs_ack_o
rlabel metal2 7682 34330 7682 34330 0 wbs_adr_i[0]
rlabel metal2 47886 35010 47886 35010 0 wbs_adr_i[10]
rlabel metal2 51382 1996 51382 1996 0 wbs_adr_i[11]
rlabel metal2 54970 35044 54970 35044 0 wbs_adr_i[12]
rlabel metal2 58466 34398 58466 34398 0 wbs_adr_i[13]
rlabel metal2 62054 26748 62054 26748 0 wbs_adr_i[14]
rlabel metal2 65550 30896 65550 30896 0 wbs_adr_i[15]
rlabel metal2 69138 1860 69138 1860 0 wbs_adr_i[16]
rlabel metal2 72634 34279 72634 34279 0 wbs_adr_i[17]
rlabel metal2 76222 33650 76222 33650 0 wbs_adr_i[18]
rlabel metal2 79718 33004 79718 33004 0 wbs_adr_i[19]
rlabel metal2 12374 32256 12374 32256 0 wbs_adr_i[1]
rlabel metal2 83306 23960 83306 23960 0 wbs_adr_i[20]
rlabel metal2 86894 33038 86894 33038 0 wbs_adr_i[21]
rlabel metal2 90390 35027 90390 35027 0 wbs_adr_i[22]
rlabel metal2 93978 34432 93978 34432 0 wbs_adr_i[23]
rlabel metal2 97474 33684 97474 33684 0 wbs_adr_i[24]
rlabel metal2 101062 33072 101062 33072 0 wbs_adr_i[25]
rlabel metal2 104558 1792 104558 1792 0 wbs_adr_i[26]
rlabel metal2 108146 2098 108146 2098 0 wbs_adr_i[27]
rlabel metal2 113850 35938 113850 35938 0 wbs_adr_i[28]
rlabel metal2 115230 33752 115230 33752 0 wbs_adr_i[29]
rlabel metal2 17066 1860 17066 1860 0 wbs_adr_i[2]
rlabel metal2 130778 72566 130778 72566 0 wbs_adr_i[30]
rlabel metal2 122314 3254 122314 3254 0 wbs_adr_i[31]
rlabel metal2 21850 33599 21850 33599 0 wbs_adr_i[3]
rlabel metal2 26542 32970 26542 32970 0 wbs_adr_i[4]
rlabel metal2 30130 34364 30130 34364 0 wbs_adr_i[5]
rlabel metal2 33626 27428 33626 27428 0 wbs_adr_i[6]
rlabel metal2 37214 1860 37214 1860 0 wbs_adr_i[7]
rlabel metal2 40710 30862 40710 30862 0 wbs_adr_i[8]
rlabel metal2 44298 31576 44298 31576 0 wbs_adr_i[9]
rlabel metal2 4094 23280 4094 23280 0 wbs_cyc_i
rlabel metal1 65320 57222 65320 57222 0 wbs_dat_i[0]
rlabel metal2 48990 32290 48990 32290 0 wbs_dat_i[10]
rlabel metal2 52578 32239 52578 32239 0 wbs_dat_i[11]
rlabel metal2 56074 31610 56074 31610 0 wbs_dat_i[12]
rlabel metal2 59662 30216 59662 30216 0 wbs_dat_i[13]
rlabel metal2 63250 30250 63250 30250 0 wbs_dat_i[14]
rlabel metal2 66746 2030 66746 2030 0 wbs_dat_i[15]
rlabel metal3 98877 58684 98877 58684 0 wbs_dat_i[16]
rlabel metal2 73830 25371 73830 25371 0 wbs_dat_i[17]
rlabel metal2 77418 28822 77418 28822 0 wbs_dat_i[18]
rlabel metal2 80914 35112 80914 35112 0 wbs_dat_i[19]
rlabel metal2 13570 26034 13570 26034 0 wbs_dat_i[1]
rlabel metal2 84502 35758 84502 35758 0 wbs_dat_i[20]
rlabel metal2 87998 30879 87998 30879 0 wbs_dat_i[21]
rlabel metal3 110055 55828 110055 55828 0 wbs_dat_i[22]
rlabel metal2 95174 22634 95174 22634 0 wbs_dat_i[23]
rlabel metal2 98670 2064 98670 2064 0 wbs_dat_i[24]
rlabel metal2 102258 31644 102258 31644 0 wbs_dat_i[25]
rlabel metal2 105754 35775 105754 35775 0 wbs_dat_i[26]
rlabel metal2 109342 30930 109342 30930 0 wbs_dat_i[27]
rlabel metal2 112838 32358 112838 32358 0 wbs_dat_i[28]
rlabel metal2 116426 35554 116426 35554 0 wbs_dat_i[29]
rlabel metal2 18262 35707 18262 35707 0 wbs_dat_i[2]
rlabel metal2 119922 1894 119922 1894 0 wbs_dat_i[30]
rlabel metal2 123273 340 123273 340 0 wbs_dat_i[31]
rlabel metal2 23046 36404 23046 36404 0 wbs_dat_i[3]
rlabel metal2 27738 1656 27738 1656 0 wbs_dat_i[4]
rlabel metal2 31326 26714 31326 26714 0 wbs_dat_i[5]
rlabel metal2 34822 33667 34822 33667 0 wbs_dat_i[6]
rlabel metal2 38410 26731 38410 26731 0 wbs_dat_i[7]
rlabel metal2 41906 35724 41906 35724 0 wbs_dat_i[8]
rlabel metal2 45494 2574 45494 2574 0 wbs_dat_i[9]
rlabel metal2 9982 30182 9982 30182 0 wbs_dat_o[0]
rlabel metal2 50186 4002 50186 4002 0 wbs_dat_o[10]
rlabel metal2 53774 23263 53774 23263 0 wbs_dat_o[11]
rlabel metal2 57270 28142 57270 28142 0 wbs_dat_o[12]
rlabel metal2 60858 33616 60858 33616 0 wbs_dat_o[13]
rlabel metal2 64354 22600 64354 22600 0 wbs_dat_o[14]
rlabel metal2 67942 32324 67942 32324 0 wbs_dat_o[15]
rlabel metal2 71530 2608 71530 2608 0 wbs_dat_o[16]
rlabel metal2 75026 24691 75026 24691 0 wbs_dat_o[17]
rlabel metal2 78614 3288 78614 3288 0 wbs_dat_o[18]
rlabel metal2 82110 20526 82110 20526 0 wbs_dat_o[19]
rlabel metal2 14766 25354 14766 25354 0 wbs_dat_o[1]
rlabel metal2 85698 6722 85698 6722 0 wbs_dat_o[20]
rlabel metal2 89194 3271 89194 3271 0 wbs_dat_o[21]
rlabel metal2 92782 23994 92782 23994 0 wbs_dat_o[22]
rlabel metal2 96278 4648 96278 4648 0 wbs_dat_o[23]
rlabel metal2 99866 24674 99866 24674 0 wbs_dat_o[24]
rlabel metal2 103362 33718 103362 33718 0 wbs_dat_o[25]
rlabel metal1 114126 57358 114126 57358 0 wbs_dat_o[26]
rlabel metal2 110538 1860 110538 1860 0 wbs_dat_o[27]
rlabel metal1 116840 58378 116840 58378 0 wbs_dat_o[28]
rlabel metal2 117622 34534 117622 34534 0 wbs_dat_o[29]
rlabel metal2 19458 5328 19458 5328 0 wbs_dat_o[2]
rlabel metal2 130962 73212 130962 73212 0 wbs_dat_o[30]
rlabel metal2 124706 1656 124706 1656 0 wbs_dat_o[31]
rlabel metal2 24242 3968 24242 3968 0 wbs_dat_o[3]
rlabel metal2 118174 43588 118174 43588 0 wbs_dat_o[4]
rlabel metal1 78108 55862 78108 55862 0 wbs_dat_o[5]
rlabel metal2 36018 8116 36018 8116 0 wbs_dat_o[6]
rlabel metal2 39606 1724 39606 1724 0 wbs_dat_o[7]
rlabel metal2 43102 8796 43102 8796 0 wbs_dat_o[8]
rlabel metal2 46690 5362 46690 5362 0 wbs_dat_o[9]
rlabel metal2 116886 45305 116886 45305 0 wbs_sel_i[0]
rlabel metal2 15962 1962 15962 1962 0 wbs_sel_i[1]
rlabel metal2 20654 12944 20654 12944 0 wbs_sel_i[2]
rlabel metal2 25346 29502 25346 29502 0 wbs_sel_i[3]
rlabel metal2 5290 2574 5290 2574 0 wbs_stb_i
rlabel metal2 6486 3254 6486 3254 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
