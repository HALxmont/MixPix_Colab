`default_nettype none

module PD_M1_M2(
    
`ifdef USE_POWER_PINS
    input   VDD,
    input   VSS,
`endif
    
    input  PD1,
    input  PD2,
    input  PD3,
    input  PD4,
    input  PD5,
    input  PD6,
    input  PD7,
    input  PD8,
    input  PD9,
    input  PD10,
    input  PD11,
    input  PD12,

);




endmodule
`default_nettype wire

