magic
tech sky130A
magscale 1 2
timestamp 1678372861
<< nwell >>
rect 8980 2610 9500 2700
rect 8960 2130 9050 2610
rect 9270 2500 9500 2610
rect 12370 -3310 12580 -3290
rect 12170 -3320 12580 -3310
rect 12400 -3490 12490 -3320
rect 12400 -3870 12510 -3490
<< pwell >>
rect -3650 4740 -3092 5310
rect -2360 4740 -1802 5310
rect -1070 4740 -512 5310
rect 220 4740 778 5310
rect 1510 4740 2068 5310
rect 2800 4740 3358 5310
rect 4090 4740 4648 5310
rect 5380 4740 5938 5310
rect 6670 4740 7228 5310
rect 7960 4740 8518 5310
rect 9250 4740 9808 5310
rect -4940 4100 -4382 4670
rect -3660 4100 -3102 4670
rect -2360 4100 -1802 4670
rect -1080 4100 -522 4670
rect 220 4100 778 4670
rect 1500 4100 2058 4670
rect 2800 4100 3358 4670
rect 4080 4100 4638 4670
rect 5380 4100 5938 4670
rect 6660 4100 7218 4670
rect 7960 4100 8518 4670
rect 9240 4100 9798 4670
<< nmoslvt >>
rect -3440 5054 -3240 5114
rect -3440 4936 -3240 4996
rect -2150 5054 -1950 5114
rect -2150 4936 -1950 4996
rect -860 5054 -660 5114
rect -860 4936 -660 4996
rect 430 5054 630 5114
rect 430 4936 630 4996
rect 1720 5054 1920 5114
rect 1720 4936 1920 4996
rect 3010 5054 3210 5114
rect 3010 4936 3210 4996
rect 4300 5054 4500 5114
rect 4300 4936 4500 4996
rect 5590 5054 5790 5114
rect 5590 4936 5790 4996
rect 6880 5054 7080 5114
rect 6880 4936 7080 4996
rect 8170 5054 8370 5114
rect 8170 4936 8370 4996
rect 9460 5054 9660 5114
rect 9460 4936 9660 4996
rect -4730 4414 -4530 4474
rect -4730 4296 -4530 4356
rect -3450 4414 -3250 4474
rect -3450 4296 -3250 4356
rect -2150 4414 -1950 4474
rect -2150 4296 -1950 4356
rect -870 4414 -670 4474
rect -870 4296 -670 4356
rect 430 4414 630 4474
rect 430 4296 630 4356
rect 1710 4414 1910 4474
rect 1710 4296 1910 4356
rect 3010 4414 3210 4474
rect 3010 4296 3210 4356
rect 4290 4414 4490 4474
rect 4290 4296 4490 4356
rect 5590 4414 5790 4474
rect 5590 4296 5790 4356
rect 6870 4414 7070 4474
rect 6870 4296 7070 4356
rect 8170 4414 8370 4474
rect 8170 4296 8370 4356
rect 9450 4414 9650 4474
rect 9450 4296 9650 4356
<< ndiff >>
rect -3440 5160 -3240 5172
rect -3440 5126 -3428 5160
rect -3252 5126 -3240 5160
rect -3440 5114 -3240 5126
rect -3440 5042 -3240 5054
rect -3440 5008 -3428 5042
rect -3252 5008 -3240 5042
rect -3440 4996 -3240 5008
rect -3440 4924 -3240 4936
rect -3440 4890 -3428 4924
rect -3252 4890 -3240 4924
rect -3440 4878 -3240 4890
rect -2150 5160 -1950 5172
rect -2150 5126 -2138 5160
rect -1962 5126 -1950 5160
rect -2150 5114 -1950 5126
rect -2150 5042 -1950 5054
rect -2150 5008 -2138 5042
rect -1962 5008 -1950 5042
rect -2150 4996 -1950 5008
rect -2150 4924 -1950 4936
rect -2150 4890 -2138 4924
rect -1962 4890 -1950 4924
rect -2150 4878 -1950 4890
rect -860 5160 -660 5172
rect -860 5126 -848 5160
rect -672 5126 -660 5160
rect -860 5114 -660 5126
rect -860 5042 -660 5054
rect -860 5008 -848 5042
rect -672 5008 -660 5042
rect -860 4996 -660 5008
rect -860 4924 -660 4936
rect -860 4890 -848 4924
rect -672 4890 -660 4924
rect -860 4878 -660 4890
rect 430 5160 630 5172
rect 430 5126 442 5160
rect 618 5126 630 5160
rect 430 5114 630 5126
rect 430 5042 630 5054
rect 430 5008 442 5042
rect 618 5008 630 5042
rect 430 4996 630 5008
rect 430 4924 630 4936
rect 430 4890 442 4924
rect 618 4890 630 4924
rect 430 4878 630 4890
rect 1720 5160 1920 5172
rect 1720 5126 1732 5160
rect 1908 5126 1920 5160
rect 1720 5114 1920 5126
rect 1720 5042 1920 5054
rect 1720 5008 1732 5042
rect 1908 5008 1920 5042
rect 1720 4996 1920 5008
rect 1720 4924 1920 4936
rect 1720 4890 1732 4924
rect 1908 4890 1920 4924
rect 1720 4878 1920 4890
rect 3010 5160 3210 5172
rect 3010 5126 3022 5160
rect 3198 5126 3210 5160
rect 3010 5114 3210 5126
rect 3010 5042 3210 5054
rect 3010 5008 3022 5042
rect 3198 5008 3210 5042
rect 3010 4996 3210 5008
rect 3010 4924 3210 4936
rect 3010 4890 3022 4924
rect 3198 4890 3210 4924
rect 3010 4878 3210 4890
rect 4300 5160 4500 5172
rect 4300 5126 4312 5160
rect 4488 5126 4500 5160
rect 4300 5114 4500 5126
rect 4300 5042 4500 5054
rect 4300 5008 4312 5042
rect 4488 5008 4500 5042
rect 4300 4996 4500 5008
rect 4300 4924 4500 4936
rect 4300 4890 4312 4924
rect 4488 4890 4500 4924
rect 4300 4878 4500 4890
rect 5590 5160 5790 5172
rect 5590 5126 5602 5160
rect 5778 5126 5790 5160
rect 5590 5114 5790 5126
rect 5590 5042 5790 5054
rect 5590 5008 5602 5042
rect 5778 5008 5790 5042
rect 5590 4996 5790 5008
rect 5590 4924 5790 4936
rect 5590 4890 5602 4924
rect 5778 4890 5790 4924
rect 5590 4878 5790 4890
rect 6880 5160 7080 5172
rect 6880 5126 6892 5160
rect 7068 5126 7080 5160
rect 6880 5114 7080 5126
rect 6880 5042 7080 5054
rect 6880 5008 6892 5042
rect 7068 5008 7080 5042
rect 6880 4996 7080 5008
rect 6880 4924 7080 4936
rect 6880 4890 6892 4924
rect 7068 4890 7080 4924
rect 6880 4878 7080 4890
rect 8170 5160 8370 5172
rect 8170 5126 8182 5160
rect 8358 5126 8370 5160
rect 8170 5114 8370 5126
rect 8170 5042 8370 5054
rect 8170 5008 8182 5042
rect 8358 5008 8370 5042
rect 8170 4996 8370 5008
rect 8170 4924 8370 4936
rect 8170 4890 8182 4924
rect 8358 4890 8370 4924
rect 8170 4878 8370 4890
rect 9460 5160 9660 5172
rect 9460 5126 9472 5160
rect 9648 5126 9660 5160
rect 9460 5114 9660 5126
rect 9460 5042 9660 5054
rect 9460 5008 9472 5042
rect 9648 5008 9660 5042
rect 9460 4996 9660 5008
rect 9460 4924 9660 4936
rect 9460 4890 9472 4924
rect 9648 4890 9660 4924
rect 9460 4878 9660 4890
rect -4730 4520 -4530 4532
rect -4730 4486 -4718 4520
rect -4542 4486 -4530 4520
rect -4730 4474 -4530 4486
rect -4730 4402 -4530 4414
rect -4730 4368 -4718 4402
rect -4542 4368 -4530 4402
rect -4730 4356 -4530 4368
rect -4730 4284 -4530 4296
rect -4730 4250 -4718 4284
rect -4542 4250 -4530 4284
rect -4730 4238 -4530 4250
rect -3450 4520 -3250 4532
rect -3450 4486 -3438 4520
rect -3262 4486 -3250 4520
rect -3450 4474 -3250 4486
rect -3450 4402 -3250 4414
rect -3450 4368 -3438 4402
rect -3262 4368 -3250 4402
rect -3450 4356 -3250 4368
rect -3450 4284 -3250 4296
rect -3450 4250 -3438 4284
rect -3262 4250 -3250 4284
rect -3450 4238 -3250 4250
rect -2150 4520 -1950 4532
rect -2150 4486 -2138 4520
rect -1962 4486 -1950 4520
rect -2150 4474 -1950 4486
rect -2150 4402 -1950 4414
rect -2150 4368 -2138 4402
rect -1962 4368 -1950 4402
rect -2150 4356 -1950 4368
rect -2150 4284 -1950 4296
rect -2150 4250 -2138 4284
rect -1962 4250 -1950 4284
rect -2150 4238 -1950 4250
rect -870 4520 -670 4532
rect -870 4486 -858 4520
rect -682 4486 -670 4520
rect -870 4474 -670 4486
rect -870 4402 -670 4414
rect -870 4368 -858 4402
rect -682 4368 -670 4402
rect -870 4356 -670 4368
rect -870 4284 -670 4296
rect -870 4250 -858 4284
rect -682 4250 -670 4284
rect -870 4238 -670 4250
rect 430 4520 630 4532
rect 430 4486 442 4520
rect 618 4486 630 4520
rect 430 4474 630 4486
rect 430 4402 630 4414
rect 430 4368 442 4402
rect 618 4368 630 4402
rect 430 4356 630 4368
rect 430 4284 630 4296
rect 430 4250 442 4284
rect 618 4250 630 4284
rect 430 4238 630 4250
rect 1710 4520 1910 4532
rect 1710 4486 1722 4520
rect 1898 4486 1910 4520
rect 1710 4474 1910 4486
rect 1710 4402 1910 4414
rect 1710 4368 1722 4402
rect 1898 4368 1910 4402
rect 1710 4356 1910 4368
rect 1710 4284 1910 4296
rect 1710 4250 1722 4284
rect 1898 4250 1910 4284
rect 1710 4238 1910 4250
rect 3010 4520 3210 4532
rect 3010 4486 3022 4520
rect 3198 4486 3210 4520
rect 3010 4474 3210 4486
rect 3010 4402 3210 4414
rect 3010 4368 3022 4402
rect 3198 4368 3210 4402
rect 3010 4356 3210 4368
rect 3010 4284 3210 4296
rect 3010 4250 3022 4284
rect 3198 4250 3210 4284
rect 3010 4238 3210 4250
rect 4290 4520 4490 4532
rect 4290 4486 4302 4520
rect 4478 4486 4490 4520
rect 4290 4474 4490 4486
rect 4290 4402 4490 4414
rect 4290 4368 4302 4402
rect 4478 4368 4490 4402
rect 4290 4356 4490 4368
rect 4290 4284 4490 4296
rect 4290 4250 4302 4284
rect 4478 4250 4490 4284
rect 4290 4238 4490 4250
rect 5590 4520 5790 4532
rect 5590 4486 5602 4520
rect 5778 4486 5790 4520
rect 5590 4474 5790 4486
rect 5590 4402 5790 4414
rect 5590 4368 5602 4402
rect 5778 4368 5790 4402
rect 5590 4356 5790 4368
rect 5590 4284 5790 4296
rect 5590 4250 5602 4284
rect 5778 4250 5790 4284
rect 5590 4238 5790 4250
rect 6870 4520 7070 4532
rect 6870 4486 6882 4520
rect 7058 4486 7070 4520
rect 6870 4474 7070 4486
rect 6870 4402 7070 4414
rect 6870 4368 6882 4402
rect 7058 4368 7070 4402
rect 6870 4356 7070 4368
rect 6870 4284 7070 4296
rect 6870 4250 6882 4284
rect 7058 4250 7070 4284
rect 6870 4238 7070 4250
rect 8170 4520 8370 4532
rect 8170 4486 8182 4520
rect 8358 4486 8370 4520
rect 8170 4474 8370 4486
rect 8170 4402 8370 4414
rect 8170 4368 8182 4402
rect 8358 4368 8370 4402
rect 8170 4356 8370 4368
rect 8170 4284 8370 4296
rect 8170 4250 8182 4284
rect 8358 4250 8370 4284
rect 8170 4238 8370 4250
rect 9450 4520 9650 4532
rect 9450 4486 9462 4520
rect 9638 4486 9650 4520
rect 9450 4474 9650 4486
rect 9450 4402 9650 4414
rect 9450 4368 9462 4402
rect 9638 4368 9650 4402
rect 9450 4356 9650 4368
rect 9450 4284 9650 4296
rect 9450 4250 9462 4284
rect 9638 4250 9650 4284
rect 9450 4238 9650 4250
<< ndiffc >>
rect -3428 5126 -3252 5160
rect -3428 5008 -3252 5042
rect -3428 4890 -3252 4924
rect -2138 5126 -1962 5160
rect -2138 5008 -1962 5042
rect -2138 4890 -1962 4924
rect -848 5126 -672 5160
rect -848 5008 -672 5042
rect -848 4890 -672 4924
rect 442 5126 618 5160
rect 442 5008 618 5042
rect 442 4890 618 4924
rect 1732 5126 1908 5160
rect 1732 5008 1908 5042
rect 1732 4890 1908 4924
rect 3022 5126 3198 5160
rect 3022 5008 3198 5042
rect 3022 4890 3198 4924
rect 4312 5126 4488 5160
rect 4312 5008 4488 5042
rect 4312 4890 4488 4924
rect 5602 5126 5778 5160
rect 5602 5008 5778 5042
rect 5602 4890 5778 4924
rect 6892 5126 7068 5160
rect 6892 5008 7068 5042
rect 6892 4890 7068 4924
rect 8182 5126 8358 5160
rect 8182 5008 8358 5042
rect 8182 4890 8358 4924
rect 9472 5126 9648 5160
rect 9472 5008 9648 5042
rect 9472 4890 9648 4924
rect -4718 4486 -4542 4520
rect -4718 4368 -4542 4402
rect -4718 4250 -4542 4284
rect -3438 4486 -3262 4520
rect -3438 4368 -3262 4402
rect -3438 4250 -3262 4284
rect -2138 4486 -1962 4520
rect -2138 4368 -1962 4402
rect -2138 4250 -1962 4284
rect -858 4486 -682 4520
rect -858 4368 -682 4402
rect -858 4250 -682 4284
rect 442 4486 618 4520
rect 442 4368 618 4402
rect 442 4250 618 4284
rect 1722 4486 1898 4520
rect 1722 4368 1898 4402
rect 1722 4250 1898 4284
rect 3022 4486 3198 4520
rect 3022 4368 3198 4402
rect 3022 4250 3198 4284
rect 4302 4486 4478 4520
rect 4302 4368 4478 4402
rect 4302 4250 4478 4284
rect 5602 4486 5778 4520
rect 5602 4368 5778 4402
rect 5602 4250 5778 4284
rect 6882 4486 7058 4520
rect 6882 4368 7058 4402
rect 6882 4250 7058 4284
rect 8182 4486 8358 4520
rect 8182 4368 8358 4402
rect 8182 4250 8358 4284
rect 9462 4486 9638 4520
rect 9462 4368 9638 4402
rect 9462 4250 9638 4284
<< psubdiff >>
rect -3614 5240 -3518 5274
rect -3224 5240 -3128 5274
rect -3614 5178 -3580 5240
rect -3162 5178 -3128 5240
rect -3614 4810 -3580 4872
rect -3162 4810 -3128 4872
rect -3614 4776 -3518 4810
rect -3224 4776 -3128 4810
rect -2324 5240 -2228 5274
rect -1934 5240 -1838 5274
rect -2324 5178 -2290 5240
rect -1872 5178 -1838 5240
rect -2324 4810 -2290 4872
rect -1872 4810 -1838 4872
rect -2324 4776 -2228 4810
rect -1934 4776 -1838 4810
rect -1034 5240 -938 5274
rect -644 5240 -548 5274
rect -1034 5178 -1000 5240
rect -582 5178 -548 5240
rect -1034 4810 -1000 4872
rect -582 4810 -548 4872
rect -1034 4776 -938 4810
rect -644 4776 -548 4810
rect 256 5240 352 5274
rect 646 5240 742 5274
rect 256 5178 290 5240
rect 708 5178 742 5240
rect 256 4810 290 4872
rect 708 4810 742 4872
rect 256 4776 352 4810
rect 646 4776 742 4810
rect 1546 5240 1642 5274
rect 1936 5240 2032 5274
rect 1546 5178 1580 5240
rect 1998 5178 2032 5240
rect 1546 4810 1580 4872
rect 1998 4810 2032 4872
rect 1546 4776 1642 4810
rect 1936 4776 2032 4810
rect 2836 5240 2932 5274
rect 3226 5240 3322 5274
rect 2836 5178 2870 5240
rect 3288 5178 3322 5240
rect 2836 4810 2870 4872
rect 3288 4810 3322 4872
rect 2836 4776 2932 4810
rect 3226 4776 3322 4810
rect 4126 5240 4222 5274
rect 4516 5240 4612 5274
rect 4126 5178 4160 5240
rect 4578 5178 4612 5240
rect 4126 4810 4160 4872
rect 4578 4810 4612 4872
rect 4126 4776 4222 4810
rect 4516 4776 4612 4810
rect 5416 5240 5512 5274
rect 5806 5240 5902 5274
rect 5416 5178 5450 5240
rect 5868 5178 5902 5240
rect 5416 4810 5450 4872
rect 5868 4810 5902 4872
rect 5416 4776 5512 4810
rect 5806 4776 5902 4810
rect 6706 5240 6802 5274
rect 7096 5240 7192 5274
rect 6706 5178 6740 5240
rect 7158 5178 7192 5240
rect 6706 4810 6740 4872
rect 7158 4810 7192 4872
rect 6706 4776 6802 4810
rect 7096 4776 7192 4810
rect 7996 5240 8092 5274
rect 8386 5240 8482 5274
rect 7996 5178 8030 5240
rect 8448 5178 8482 5240
rect 7996 4810 8030 4872
rect 8448 4810 8482 4872
rect 7996 4776 8092 4810
rect 8386 4776 8482 4810
rect 9286 5240 9382 5274
rect 9676 5240 9772 5274
rect 9286 5178 9320 5240
rect 9738 5178 9772 5240
rect 9286 4810 9320 4872
rect 9738 4810 9772 4872
rect 9286 4776 9382 4810
rect 9676 4776 9772 4810
rect -4904 4600 -4808 4634
rect -4514 4600 -4418 4634
rect -4904 4538 -4870 4600
rect -4452 4538 -4418 4600
rect -4904 4170 -4870 4232
rect -4452 4170 -4418 4232
rect -4904 4136 -4808 4170
rect -4514 4136 -4418 4170
rect -3624 4600 -3528 4634
rect -3234 4600 -3138 4634
rect -3624 4538 -3590 4600
rect -3172 4538 -3138 4600
rect -3624 4170 -3590 4232
rect -3172 4170 -3138 4232
rect -3624 4136 -3528 4170
rect -3234 4136 -3138 4170
rect -2324 4600 -2228 4634
rect -1934 4600 -1838 4634
rect -2324 4538 -2290 4600
rect -1872 4538 -1838 4600
rect -2324 4170 -2290 4232
rect -1872 4170 -1838 4232
rect -2324 4136 -2228 4170
rect -1934 4136 -1838 4170
rect -1044 4600 -948 4634
rect -654 4600 -558 4634
rect -1044 4538 -1010 4600
rect -592 4538 -558 4600
rect -1044 4170 -1010 4232
rect -592 4170 -558 4232
rect -1044 4136 -948 4170
rect -654 4136 -558 4170
rect 256 4600 352 4634
rect 646 4600 742 4634
rect 256 4538 290 4600
rect 708 4538 742 4600
rect 256 4170 290 4232
rect 708 4170 742 4232
rect 256 4136 352 4170
rect 646 4136 742 4170
rect 1536 4600 1632 4634
rect 1926 4600 2022 4634
rect 1536 4538 1570 4600
rect 1988 4538 2022 4600
rect 1536 4170 1570 4232
rect 1988 4170 2022 4232
rect 1536 4136 1632 4170
rect 1926 4136 2022 4170
rect 2836 4600 2932 4634
rect 3226 4600 3322 4634
rect 2836 4538 2870 4600
rect 3288 4538 3322 4600
rect 2836 4170 2870 4232
rect 3288 4170 3322 4232
rect 2836 4136 2932 4170
rect 3226 4136 3322 4170
rect 4116 4600 4212 4634
rect 4506 4600 4602 4634
rect 4116 4538 4150 4600
rect 4568 4538 4602 4600
rect 4116 4170 4150 4232
rect 4568 4170 4602 4232
rect 4116 4136 4212 4170
rect 4506 4136 4602 4170
rect 5416 4600 5512 4634
rect 5806 4600 5902 4634
rect 5416 4538 5450 4600
rect 5868 4538 5902 4600
rect 5416 4170 5450 4232
rect 5868 4170 5902 4232
rect 5416 4136 5512 4170
rect 5806 4136 5902 4170
rect 6696 4600 6792 4634
rect 7086 4600 7182 4634
rect 6696 4538 6730 4600
rect 7148 4538 7182 4600
rect 6696 4170 6730 4232
rect 7148 4170 7182 4232
rect 6696 4136 6792 4170
rect 7086 4136 7182 4170
rect 7996 4600 8092 4634
rect 8386 4600 8482 4634
rect 7996 4538 8030 4600
rect 8448 4538 8482 4600
rect 7996 4170 8030 4232
rect 8448 4170 8482 4232
rect 7996 4136 8092 4170
rect 8386 4136 8482 4170
rect 9276 4600 9372 4634
rect 9666 4600 9762 4634
rect 9276 4538 9310 4600
rect 9728 4538 9762 4600
rect 9276 4170 9310 4232
rect 9728 4170 9762 4232
rect 9276 4136 9372 4170
rect 9666 4136 9762 4170
<< psubdiffcont >>
rect -3518 5240 -3224 5274
rect -3614 4872 -3580 5178
rect -3162 4872 -3128 5178
rect -3518 4776 -3224 4810
rect -2228 5240 -1934 5274
rect -2324 4872 -2290 5178
rect -1872 4872 -1838 5178
rect -2228 4776 -1934 4810
rect -938 5240 -644 5274
rect -1034 4872 -1000 5178
rect -582 4872 -548 5178
rect -938 4776 -644 4810
rect 352 5240 646 5274
rect 256 4872 290 5178
rect 708 4872 742 5178
rect 352 4776 646 4810
rect 1642 5240 1936 5274
rect 1546 4872 1580 5178
rect 1998 4872 2032 5178
rect 1642 4776 1936 4810
rect 2932 5240 3226 5274
rect 2836 4872 2870 5178
rect 3288 4872 3322 5178
rect 2932 4776 3226 4810
rect 4222 5240 4516 5274
rect 4126 4872 4160 5178
rect 4578 4872 4612 5178
rect 4222 4776 4516 4810
rect 5512 5240 5806 5274
rect 5416 4872 5450 5178
rect 5868 4872 5902 5178
rect 5512 4776 5806 4810
rect 6802 5240 7096 5274
rect 6706 4872 6740 5178
rect 7158 4872 7192 5178
rect 6802 4776 7096 4810
rect 8092 5240 8386 5274
rect 7996 4872 8030 5178
rect 8448 4872 8482 5178
rect 8092 4776 8386 4810
rect 9382 5240 9676 5274
rect 9286 4872 9320 5178
rect 9738 4872 9772 5178
rect 9382 4776 9676 4810
rect -4808 4600 -4514 4634
rect -4904 4232 -4870 4538
rect -4452 4232 -4418 4538
rect -4808 4136 -4514 4170
rect -3528 4600 -3234 4634
rect -3624 4232 -3590 4538
rect -3172 4232 -3138 4538
rect -3528 4136 -3234 4170
rect -2228 4600 -1934 4634
rect -2324 4232 -2290 4538
rect -1872 4232 -1838 4538
rect -2228 4136 -1934 4170
rect -948 4600 -654 4634
rect -1044 4232 -1010 4538
rect -592 4232 -558 4538
rect -948 4136 -654 4170
rect 352 4600 646 4634
rect 256 4232 290 4538
rect 708 4232 742 4538
rect 352 4136 646 4170
rect 1632 4600 1926 4634
rect 1536 4232 1570 4538
rect 1988 4232 2022 4538
rect 1632 4136 1926 4170
rect 2932 4600 3226 4634
rect 2836 4232 2870 4538
rect 3288 4232 3322 4538
rect 2932 4136 3226 4170
rect 4212 4600 4506 4634
rect 4116 4232 4150 4538
rect 4568 4232 4602 4538
rect 4212 4136 4506 4170
rect 5512 4600 5806 4634
rect 5416 4232 5450 4538
rect 5868 4232 5902 4538
rect 5512 4136 5806 4170
rect 6792 4600 7086 4634
rect 6696 4232 6730 4538
rect 7148 4232 7182 4538
rect 6792 4136 7086 4170
rect 8092 4600 8386 4634
rect 7996 4232 8030 4538
rect 8448 4232 8482 4538
rect 8092 4136 8386 4170
rect 9372 4600 9666 4634
rect 9276 4232 9310 4538
rect 9728 4232 9762 4538
rect 9372 4136 9666 4170
<< poly >>
rect -3528 5114 -3462 5117
rect -3528 5101 -3440 5114
rect -3528 5067 -3512 5101
rect -3478 5067 -3440 5101
rect -3528 5054 -3440 5067
rect -3240 5054 -3214 5114
rect -3528 5051 -3462 5054
rect -3528 4996 -3462 4999
rect -3528 4983 -3440 4996
rect -3528 4949 -3512 4983
rect -3478 4949 -3440 4983
rect -3528 4936 -3440 4949
rect -3240 4936 -3214 4996
rect -3528 4933 -3462 4936
rect -2238 5114 -2172 5117
rect -2238 5101 -2150 5114
rect -2238 5067 -2222 5101
rect -2188 5067 -2150 5101
rect -2238 5054 -2150 5067
rect -1950 5054 -1924 5114
rect -2238 5051 -2172 5054
rect -2238 4996 -2172 4999
rect -2238 4983 -2150 4996
rect -2238 4949 -2222 4983
rect -2188 4949 -2150 4983
rect -2238 4936 -2150 4949
rect -1950 4936 -1924 4996
rect -2238 4933 -2172 4936
rect -948 5114 -882 5117
rect -948 5101 -860 5114
rect -948 5067 -932 5101
rect -898 5067 -860 5101
rect -948 5054 -860 5067
rect -660 5054 -634 5114
rect -948 5051 -882 5054
rect -948 4996 -882 4999
rect -948 4983 -860 4996
rect -948 4949 -932 4983
rect -898 4949 -860 4983
rect -948 4936 -860 4949
rect -660 4936 -634 4996
rect -948 4933 -882 4936
rect 342 5114 408 5117
rect 342 5101 430 5114
rect 342 5067 358 5101
rect 392 5067 430 5101
rect 342 5054 430 5067
rect 630 5054 656 5114
rect 342 5051 408 5054
rect 342 4996 408 4999
rect 342 4983 430 4996
rect 342 4949 358 4983
rect 392 4949 430 4983
rect 342 4936 430 4949
rect 630 4936 656 4996
rect 342 4933 408 4936
rect 1632 5114 1698 5117
rect 1632 5101 1720 5114
rect 1632 5067 1648 5101
rect 1682 5067 1720 5101
rect 1632 5054 1720 5067
rect 1920 5054 1946 5114
rect 1632 5051 1698 5054
rect 1632 4996 1698 4999
rect 1632 4983 1720 4996
rect 1632 4949 1648 4983
rect 1682 4949 1720 4983
rect 1632 4936 1720 4949
rect 1920 4936 1946 4996
rect 1632 4933 1698 4936
rect 2922 5114 2988 5117
rect 2922 5101 3010 5114
rect 2922 5067 2938 5101
rect 2972 5067 3010 5101
rect 2922 5054 3010 5067
rect 3210 5054 3236 5114
rect 2922 5051 2988 5054
rect 2922 4996 2988 4999
rect 2922 4983 3010 4996
rect 2922 4949 2938 4983
rect 2972 4949 3010 4983
rect 2922 4936 3010 4949
rect 3210 4936 3236 4996
rect 2922 4933 2988 4936
rect 4212 5114 4278 5117
rect 4212 5101 4300 5114
rect 4212 5067 4228 5101
rect 4262 5067 4300 5101
rect 4212 5054 4300 5067
rect 4500 5054 4526 5114
rect 4212 5051 4278 5054
rect 4212 4996 4278 4999
rect 4212 4983 4300 4996
rect 4212 4949 4228 4983
rect 4262 4949 4300 4983
rect 4212 4936 4300 4949
rect 4500 4936 4526 4996
rect 4212 4933 4278 4936
rect 5502 5114 5568 5117
rect 5502 5101 5590 5114
rect 5502 5067 5518 5101
rect 5552 5067 5590 5101
rect 5502 5054 5590 5067
rect 5790 5054 5816 5114
rect 5502 5051 5568 5054
rect 5502 4996 5568 4999
rect 5502 4983 5590 4996
rect 5502 4949 5518 4983
rect 5552 4949 5590 4983
rect 5502 4936 5590 4949
rect 5790 4936 5816 4996
rect 5502 4933 5568 4936
rect 6792 5114 6858 5117
rect 6792 5101 6880 5114
rect 6792 5067 6808 5101
rect 6842 5067 6880 5101
rect 6792 5054 6880 5067
rect 7080 5054 7106 5114
rect 6792 5051 6858 5054
rect 6792 4996 6858 4999
rect 6792 4983 6880 4996
rect 6792 4949 6808 4983
rect 6842 4949 6880 4983
rect 6792 4936 6880 4949
rect 7080 4936 7106 4996
rect 6792 4933 6858 4936
rect 8082 5114 8148 5117
rect 8082 5101 8170 5114
rect 8082 5067 8098 5101
rect 8132 5067 8170 5101
rect 8082 5054 8170 5067
rect 8370 5054 8396 5114
rect 8082 5051 8148 5054
rect 8082 4996 8148 4999
rect 8082 4983 8170 4996
rect 8082 4949 8098 4983
rect 8132 4949 8170 4983
rect 8082 4936 8170 4949
rect 8370 4936 8396 4996
rect 8082 4933 8148 4936
rect 9372 5114 9438 5117
rect 9372 5101 9460 5114
rect 9372 5067 9388 5101
rect 9422 5067 9460 5101
rect 9372 5054 9460 5067
rect 9660 5054 9686 5114
rect 9372 5051 9438 5054
rect 9372 4996 9438 4999
rect 9372 4983 9460 4996
rect 9372 4949 9388 4983
rect 9422 4949 9460 4983
rect 9372 4936 9460 4949
rect 9660 4936 9686 4996
rect 9372 4933 9438 4936
rect -4818 4474 -4752 4477
rect -4818 4461 -4730 4474
rect -4818 4427 -4802 4461
rect -4768 4427 -4730 4461
rect -4818 4414 -4730 4427
rect -4530 4414 -4504 4474
rect -4818 4411 -4752 4414
rect -4818 4356 -4752 4359
rect -4818 4343 -4730 4356
rect -4818 4309 -4802 4343
rect -4768 4309 -4730 4343
rect -4818 4296 -4730 4309
rect -4530 4296 -4504 4356
rect -4818 4293 -4752 4296
rect -3538 4474 -3472 4477
rect -3538 4461 -3450 4474
rect -3538 4427 -3522 4461
rect -3488 4427 -3450 4461
rect -3538 4414 -3450 4427
rect -3250 4414 -3224 4474
rect -3538 4411 -3472 4414
rect -3538 4356 -3472 4359
rect -3538 4343 -3450 4356
rect -3538 4309 -3522 4343
rect -3488 4309 -3450 4343
rect -3538 4296 -3450 4309
rect -3250 4296 -3224 4356
rect -3538 4293 -3472 4296
rect -2238 4474 -2172 4477
rect -2238 4461 -2150 4474
rect -2238 4427 -2222 4461
rect -2188 4427 -2150 4461
rect -2238 4414 -2150 4427
rect -1950 4414 -1924 4474
rect -2238 4411 -2172 4414
rect -2238 4356 -2172 4359
rect -2238 4343 -2150 4356
rect -2238 4309 -2222 4343
rect -2188 4309 -2150 4343
rect -2238 4296 -2150 4309
rect -1950 4296 -1924 4356
rect -2238 4293 -2172 4296
rect -958 4474 -892 4477
rect -958 4461 -870 4474
rect -958 4427 -942 4461
rect -908 4427 -870 4461
rect -958 4414 -870 4427
rect -670 4414 -644 4474
rect -958 4411 -892 4414
rect -958 4356 -892 4359
rect -958 4343 -870 4356
rect -958 4309 -942 4343
rect -908 4309 -870 4343
rect -958 4296 -870 4309
rect -670 4296 -644 4356
rect -958 4293 -892 4296
rect 342 4474 408 4477
rect 342 4461 430 4474
rect 342 4427 358 4461
rect 392 4427 430 4461
rect 342 4414 430 4427
rect 630 4414 656 4474
rect 342 4411 408 4414
rect 342 4356 408 4359
rect 342 4343 430 4356
rect 342 4309 358 4343
rect 392 4309 430 4343
rect 342 4296 430 4309
rect 630 4296 656 4356
rect 342 4293 408 4296
rect 1622 4474 1688 4477
rect 1622 4461 1710 4474
rect 1622 4427 1638 4461
rect 1672 4427 1710 4461
rect 1622 4414 1710 4427
rect 1910 4414 1936 4474
rect 1622 4411 1688 4414
rect 1622 4356 1688 4359
rect 1622 4343 1710 4356
rect 1622 4309 1638 4343
rect 1672 4309 1710 4343
rect 1622 4296 1710 4309
rect 1910 4296 1936 4356
rect 1622 4293 1688 4296
rect 2922 4474 2988 4477
rect 2922 4461 3010 4474
rect 2922 4427 2938 4461
rect 2972 4427 3010 4461
rect 2922 4414 3010 4427
rect 3210 4414 3236 4474
rect 2922 4411 2988 4414
rect 2922 4356 2988 4359
rect 2922 4343 3010 4356
rect 2922 4309 2938 4343
rect 2972 4309 3010 4343
rect 2922 4296 3010 4309
rect 3210 4296 3236 4356
rect 2922 4293 2988 4296
rect 4202 4474 4268 4477
rect 4202 4461 4290 4474
rect 4202 4427 4218 4461
rect 4252 4427 4290 4461
rect 4202 4414 4290 4427
rect 4490 4414 4516 4474
rect 4202 4411 4268 4414
rect 4202 4356 4268 4359
rect 4202 4343 4290 4356
rect 4202 4309 4218 4343
rect 4252 4309 4290 4343
rect 4202 4296 4290 4309
rect 4490 4296 4516 4356
rect 4202 4293 4268 4296
rect 5502 4474 5568 4477
rect 5502 4461 5590 4474
rect 5502 4427 5518 4461
rect 5552 4427 5590 4461
rect 5502 4414 5590 4427
rect 5790 4414 5816 4474
rect 5502 4411 5568 4414
rect 5502 4356 5568 4359
rect 5502 4343 5590 4356
rect 5502 4309 5518 4343
rect 5552 4309 5590 4343
rect 5502 4296 5590 4309
rect 5790 4296 5816 4356
rect 5502 4293 5568 4296
rect 6782 4474 6848 4477
rect 6782 4461 6870 4474
rect 6782 4427 6798 4461
rect 6832 4427 6870 4461
rect 6782 4414 6870 4427
rect 7070 4414 7096 4474
rect 6782 4411 6848 4414
rect 6782 4356 6848 4359
rect 6782 4343 6870 4356
rect 6782 4309 6798 4343
rect 6832 4309 6870 4343
rect 6782 4296 6870 4309
rect 7070 4296 7096 4356
rect 6782 4293 6848 4296
rect 8082 4474 8148 4477
rect 8082 4461 8170 4474
rect 8082 4427 8098 4461
rect 8132 4427 8170 4461
rect 8082 4414 8170 4427
rect 8370 4414 8396 4474
rect 8082 4411 8148 4414
rect 8082 4356 8148 4359
rect 8082 4343 8170 4356
rect 8082 4309 8098 4343
rect 8132 4309 8170 4343
rect 8082 4296 8170 4309
rect 8370 4296 8396 4356
rect 8082 4293 8148 4296
rect 9362 4474 9428 4477
rect 9362 4461 9450 4474
rect 9362 4427 9378 4461
rect 9412 4427 9450 4461
rect 9362 4414 9450 4427
rect 9650 4414 9676 4474
rect 9362 4411 9428 4414
rect 9362 4356 9428 4359
rect 9362 4343 9450 4356
rect 9362 4309 9378 4343
rect 9412 4309 9450 4343
rect 9362 4296 9450 4309
rect 9650 4296 9676 4356
rect 9362 4293 9428 4296
<< polycont >>
rect -3512 5067 -3478 5101
rect -3512 4949 -3478 4983
rect -2222 5067 -2188 5101
rect -2222 4949 -2188 4983
rect -932 5067 -898 5101
rect -932 4949 -898 4983
rect 358 5067 392 5101
rect 358 4949 392 4983
rect 1648 5067 1682 5101
rect 1648 4949 1682 4983
rect 2938 5067 2972 5101
rect 2938 4949 2972 4983
rect 4228 5067 4262 5101
rect 4228 4949 4262 4983
rect 5518 5067 5552 5101
rect 5518 4949 5552 4983
rect 6808 5067 6842 5101
rect 6808 4949 6842 4983
rect 8098 5067 8132 5101
rect 8098 4949 8132 4983
rect 9388 5067 9422 5101
rect 9388 4949 9422 4983
rect -4802 4427 -4768 4461
rect -4802 4309 -4768 4343
rect -3522 4427 -3488 4461
rect -3522 4309 -3488 4343
rect -2222 4427 -2188 4461
rect -2222 4309 -2188 4343
rect -942 4427 -908 4461
rect -942 4309 -908 4343
rect 358 4427 392 4461
rect 358 4309 392 4343
rect 1638 4427 1672 4461
rect 1638 4309 1672 4343
rect 2938 4427 2972 4461
rect 2938 4309 2972 4343
rect 4218 4427 4252 4461
rect 4218 4309 4252 4343
rect 5518 4427 5552 4461
rect 5518 4309 5552 4343
rect 6798 4427 6832 4461
rect 6798 4309 6832 4343
rect 8098 4427 8132 4461
rect 8098 4309 8132 4343
rect 9378 4427 9412 4461
rect 9378 4309 9412 4343
<< locali >>
rect -3614 5240 -3518 5274
rect -3224 5240 -3128 5274
rect -4360 5180 -4300 5200
rect -4360 5130 -4350 5180
rect -4310 5130 -4300 5180
rect -4830 5100 -4770 5130
rect -4360 5110 -4300 5130
rect -4830 4960 -4820 5100
rect -4780 4960 -4770 5100
rect -4830 4930 -4770 4960
rect -4340 4950 -4300 5110
rect -3614 5178 -3580 5240
rect -4350 4930 -4290 4950
rect -4350 4880 -4340 4930
rect -4300 4880 -4290 4930
rect -4350 4860 -4290 4880
rect -3162 5178 -3128 5240
rect -2324 5240 -2228 5274
rect -1934 5240 -1838 5274
rect -3540 5117 -3480 5130
rect -3444 5126 -3428 5160
rect -3252 5126 -3236 5160
rect -3540 5101 -3478 5117
rect -3540 5100 -3512 5101
rect -3540 4960 -3530 5100
rect -3490 5051 -3478 5067
rect -3490 4999 -3480 5051
rect -3444 5008 -3428 5042
rect -3252 5008 -3236 5042
rect -3490 4983 -3478 4999
rect -3540 4949 -3512 4960
rect -3540 4933 -3478 4949
rect -3540 4930 -3480 4933
rect -3444 4890 -3428 4924
rect -3252 4890 -3236 4924
rect -3614 4820 -3580 4872
rect -3070 5180 -3010 5200
rect -3070 5130 -3060 5180
rect -3020 5130 -3010 5180
rect -3070 5110 -3010 5130
rect -3050 4950 -3010 5110
rect -2324 5178 -2290 5240
rect -3162 4820 -3128 4872
rect -3060 4930 -3000 4950
rect -3060 4880 -3050 4930
rect -3010 4880 -3000 4930
rect -3060 4860 -3000 4880
rect -1872 5178 -1838 5240
rect -1034 5240 -938 5274
rect -644 5240 -548 5274
rect -2250 5117 -2190 5130
rect -2154 5126 -2138 5160
rect -1962 5126 -1946 5160
rect -2250 5101 -2188 5117
rect -2250 5100 -2222 5101
rect -2250 4960 -2240 5100
rect -2200 5051 -2188 5067
rect -2200 4999 -2190 5051
rect -2154 5008 -2138 5042
rect -1962 5008 -1946 5042
rect -2200 4983 -2188 4999
rect -2250 4949 -2222 4960
rect -2250 4933 -2188 4949
rect -2250 4930 -2190 4933
rect -2154 4890 -2138 4924
rect -1962 4890 -1946 4924
rect -2324 4820 -2290 4872
rect -1780 5180 -1720 5200
rect -1780 5130 -1770 5180
rect -1730 5130 -1720 5180
rect -1780 5110 -1720 5130
rect -1760 4950 -1720 5110
rect -1034 5178 -1000 5240
rect -1872 4820 -1838 4872
rect -1770 4930 -1710 4950
rect -1770 4880 -1760 4930
rect -1720 4880 -1710 4930
rect -1770 4860 -1710 4880
rect -582 5178 -548 5240
rect 256 5240 352 5274
rect 646 5240 742 5274
rect -960 5117 -900 5130
rect -864 5126 -848 5160
rect -672 5126 -656 5160
rect -960 5101 -898 5117
rect -960 5100 -932 5101
rect -960 4960 -950 5100
rect -910 5051 -898 5067
rect -910 4999 -900 5051
rect -864 5008 -848 5042
rect -672 5008 -656 5042
rect -910 4983 -898 4999
rect -960 4949 -932 4960
rect -960 4933 -898 4949
rect -960 4930 -900 4933
rect -864 4890 -848 4924
rect -672 4890 -656 4924
rect -1034 4820 -1000 4872
rect -490 5180 -430 5200
rect -490 5130 -480 5180
rect -440 5130 -430 5180
rect -490 5110 -430 5130
rect -470 4950 -430 5110
rect 256 5178 290 5240
rect -582 4820 -548 4872
rect -480 4930 -420 4950
rect -480 4880 -470 4930
rect -430 4880 -420 4930
rect -480 4860 -420 4880
rect 708 5178 742 5240
rect 1546 5240 1642 5274
rect 1936 5240 2032 5274
rect 330 5117 390 5130
rect 426 5126 442 5160
rect 618 5126 634 5160
rect 330 5101 392 5117
rect 330 5100 358 5101
rect 330 4960 340 5100
rect 380 5051 392 5067
rect 380 4999 390 5051
rect 426 5008 442 5042
rect 618 5008 634 5042
rect 380 4983 392 4999
rect 330 4949 358 4960
rect 330 4933 392 4949
rect 330 4930 390 4933
rect 426 4890 442 4924
rect 618 4890 634 4924
rect 256 4820 290 4872
rect 800 5180 860 5200
rect 800 5130 810 5180
rect 850 5130 860 5180
rect 800 5110 860 5130
rect 820 4950 860 5110
rect 1546 5178 1580 5240
rect 708 4820 742 4872
rect 810 4930 870 4950
rect 810 4880 820 4930
rect 860 4880 870 4930
rect 810 4860 870 4880
rect 1998 5178 2032 5240
rect 2836 5240 2932 5274
rect 3226 5240 3322 5274
rect 1620 5117 1680 5130
rect 1716 5126 1732 5160
rect 1908 5126 1924 5160
rect 1620 5101 1682 5117
rect 1620 5100 1648 5101
rect 1620 4960 1630 5100
rect 1670 5051 1682 5067
rect 1670 4999 1680 5051
rect 1716 5008 1732 5042
rect 1908 5008 1924 5042
rect 1670 4983 1682 4999
rect 1620 4949 1648 4960
rect 1620 4933 1682 4949
rect 1620 4930 1680 4933
rect 1716 4890 1732 4924
rect 1908 4890 1924 4924
rect 1546 4820 1580 4872
rect 2090 5180 2150 5200
rect 2090 5130 2100 5180
rect 2140 5130 2150 5180
rect 2090 5110 2150 5130
rect 2110 4950 2150 5110
rect 2836 5178 2870 5240
rect 1998 4820 2032 4872
rect 2100 4930 2160 4950
rect 2100 4880 2110 4930
rect 2150 4880 2160 4930
rect 2100 4860 2160 4880
rect 3288 5178 3322 5240
rect 4126 5240 4222 5274
rect 4516 5240 4612 5274
rect 2910 5117 2970 5130
rect 3006 5126 3022 5160
rect 3198 5126 3214 5160
rect 2910 5101 2972 5117
rect 2910 5100 2938 5101
rect 2910 4960 2920 5100
rect 2960 5051 2972 5067
rect 2960 4999 2970 5051
rect 3006 5008 3022 5042
rect 3198 5008 3214 5042
rect 2960 4983 2972 4999
rect 2910 4949 2938 4960
rect 2910 4933 2972 4949
rect 2910 4930 2970 4933
rect 3006 4890 3022 4924
rect 3198 4890 3214 4924
rect 2836 4820 2870 4872
rect 3380 5180 3440 5200
rect 3380 5130 3390 5180
rect 3430 5130 3440 5180
rect 3380 5110 3440 5130
rect 3400 4950 3440 5110
rect 4126 5178 4160 5240
rect 3288 4820 3322 4872
rect 3390 4930 3450 4950
rect 3390 4880 3400 4930
rect 3440 4880 3450 4930
rect 3390 4860 3450 4880
rect 4578 5178 4612 5240
rect 5416 5240 5512 5274
rect 5806 5240 5902 5274
rect 4200 5117 4260 5130
rect 4296 5126 4312 5160
rect 4488 5126 4504 5160
rect 4200 5101 4262 5117
rect 4200 5100 4228 5101
rect 4200 4960 4210 5100
rect 4250 5051 4262 5067
rect 4250 4999 4260 5051
rect 4296 5008 4312 5042
rect 4488 5008 4504 5042
rect 4250 4983 4262 4999
rect 4200 4949 4228 4960
rect 4200 4933 4262 4949
rect 4200 4930 4260 4933
rect 4296 4890 4312 4924
rect 4488 4890 4504 4924
rect 4126 4820 4160 4872
rect 4670 5180 4730 5200
rect 4670 5130 4680 5180
rect 4720 5130 4730 5180
rect 4670 5110 4730 5130
rect 4690 4950 4730 5110
rect 5416 5178 5450 5240
rect 4578 4820 4612 4872
rect 4680 4930 4740 4950
rect 4680 4880 4690 4930
rect 4730 4880 4740 4930
rect 4680 4860 4740 4880
rect 5868 5178 5902 5240
rect 6706 5240 6802 5274
rect 7096 5240 7192 5274
rect 5490 5117 5550 5130
rect 5586 5126 5602 5160
rect 5778 5126 5794 5160
rect 5490 5101 5552 5117
rect 5490 5100 5518 5101
rect 5490 4960 5500 5100
rect 5540 5051 5552 5067
rect 5540 4999 5550 5051
rect 5586 5008 5602 5042
rect 5778 5008 5794 5042
rect 5540 4983 5552 4999
rect 5490 4949 5518 4960
rect 5490 4933 5552 4949
rect 5490 4930 5550 4933
rect 5586 4890 5602 4924
rect 5778 4890 5794 4924
rect 5416 4820 5450 4872
rect 5960 5180 6020 5200
rect 5960 5130 5970 5180
rect 6010 5130 6020 5180
rect 5960 5110 6020 5130
rect 5980 4950 6020 5110
rect 6706 5178 6740 5240
rect 5868 4820 5902 4872
rect 5970 4930 6030 4950
rect 5970 4880 5980 4930
rect 6020 4880 6030 4930
rect 5970 4860 6030 4880
rect 7158 5178 7192 5240
rect 7996 5240 8092 5274
rect 8386 5240 8482 5274
rect 6780 5117 6840 5130
rect 6876 5126 6892 5160
rect 7068 5126 7084 5160
rect 6780 5101 6842 5117
rect 6780 5100 6808 5101
rect 6780 4960 6790 5100
rect 6830 5051 6842 5067
rect 6830 4999 6840 5051
rect 6876 5008 6892 5042
rect 7068 5008 7084 5042
rect 6830 4983 6842 4999
rect 6780 4949 6808 4960
rect 6780 4933 6842 4949
rect 6780 4930 6840 4933
rect 6876 4890 6892 4924
rect 7068 4890 7084 4924
rect 6706 4820 6740 4872
rect 7250 5180 7310 5200
rect 7250 5130 7260 5180
rect 7300 5130 7310 5180
rect 7250 5110 7310 5130
rect 7270 4950 7310 5110
rect 7996 5178 8030 5240
rect 7158 4820 7192 4872
rect 7260 4930 7320 4950
rect 7260 4880 7270 4930
rect 7310 4880 7320 4930
rect 7260 4860 7320 4880
rect 8448 5178 8482 5240
rect 9286 5240 9382 5274
rect 9676 5240 9772 5274
rect 8070 5117 8130 5130
rect 8166 5126 8182 5160
rect 8358 5126 8374 5160
rect 8070 5101 8132 5117
rect 8070 5100 8098 5101
rect 8070 4960 8080 5100
rect 8120 5051 8132 5067
rect 8120 4999 8130 5051
rect 8166 5008 8182 5042
rect 8358 5008 8374 5042
rect 8120 4983 8132 4999
rect 8070 4949 8098 4960
rect 8070 4933 8132 4949
rect 8070 4930 8130 4933
rect 8166 4890 8182 4924
rect 8358 4890 8374 4924
rect 7996 4820 8030 4872
rect 8540 5180 8600 5200
rect 8540 5130 8550 5180
rect 8590 5130 8600 5180
rect 8540 5110 8600 5130
rect 8560 4950 8600 5110
rect 9286 5178 9320 5240
rect 8448 4820 8482 4872
rect 8550 4930 8610 4950
rect 8550 4880 8560 4930
rect 8600 4880 8610 4930
rect 8550 4860 8610 4880
rect 9738 5178 9772 5240
rect 9360 5117 9420 5130
rect 9456 5126 9472 5160
rect 9648 5126 9664 5160
rect 9360 5101 9422 5117
rect 9360 5100 9388 5101
rect 9360 4960 9370 5100
rect 9410 5051 9422 5067
rect 9410 4999 9420 5051
rect 9456 5008 9472 5042
rect 9648 5008 9664 5042
rect 9410 4983 9422 4999
rect 9360 4949 9388 4960
rect 9360 4933 9422 4949
rect 9360 4930 9420 4933
rect 9456 4890 9472 4924
rect 9648 4890 9664 4924
rect 9286 4820 9320 4872
rect 9830 5180 9890 5200
rect 9830 5130 9840 5180
rect 9880 5130 9890 5180
rect 9830 5110 9890 5130
rect 9850 4950 9890 5110
rect 9738 4820 9772 4872
rect 9840 4930 9900 4950
rect 9840 4880 9850 4930
rect 9890 4880 9900 4930
rect 9840 4860 9900 4880
rect -4940 4810 9820 4820
rect -4940 4776 -3518 4810
rect -3224 4776 -2228 4810
rect -1934 4776 -938 4810
rect -644 4776 352 4810
rect 646 4776 1642 4810
rect 1936 4776 2932 4810
rect 3226 4776 4222 4810
rect 4516 4776 5512 4810
rect 5806 4776 6802 4810
rect 7096 4776 8092 4810
rect 8386 4776 9382 4810
rect 9676 4776 9820 4810
rect -4940 4740 9820 4776
rect -4940 4634 -4880 4740
rect -4940 4600 -4808 4634
rect -4514 4600 -4418 4634
rect -4940 4538 -4870 4600
rect -4940 4232 -4904 4538
rect -4452 4538 -4418 4600
rect -4830 4477 -4770 4490
rect -4734 4486 -4718 4520
rect -4542 4486 -4526 4520
rect -4830 4461 -4768 4477
rect -4830 4460 -4802 4461
rect -4830 4320 -4820 4460
rect -4780 4411 -4768 4427
rect -4780 4359 -4770 4411
rect -4734 4368 -4718 4402
rect -4542 4368 -4526 4402
rect -4780 4343 -4768 4359
rect -4830 4309 -4802 4320
rect -4830 4293 -4768 4309
rect -4830 4290 -4770 4293
rect -4734 4250 -4718 4284
rect -4542 4250 -4526 4284
rect -4940 4180 -4870 4232
rect -4452 4180 -4418 4232
rect -3624 4600 -3528 4634
rect -3234 4600 -3138 4634
rect -3624 4538 -3590 4600
rect -3172 4538 -3138 4600
rect -3550 4477 -3490 4490
rect -3454 4486 -3438 4520
rect -3262 4486 -3246 4520
rect -3550 4461 -3488 4477
rect -3550 4460 -3522 4461
rect -3550 4320 -3540 4460
rect -3500 4411 -3488 4427
rect -3500 4359 -3490 4411
rect -3454 4368 -3438 4402
rect -3262 4368 -3246 4402
rect -3500 4343 -3488 4359
rect -3550 4309 -3522 4320
rect -3550 4293 -3488 4309
rect -3550 4290 -3490 4293
rect -3454 4250 -3438 4284
rect -3262 4250 -3246 4284
rect -3624 4180 -3590 4232
rect -3172 4180 -3138 4232
rect -2324 4600 -2228 4634
rect -1934 4600 -1838 4634
rect -2324 4538 -2290 4600
rect -1872 4538 -1838 4600
rect -2250 4477 -2190 4490
rect -2154 4486 -2138 4520
rect -1962 4486 -1946 4520
rect -2250 4461 -2188 4477
rect -2250 4460 -2222 4461
rect -2250 4320 -2240 4460
rect -2200 4411 -2188 4427
rect -2200 4359 -2190 4411
rect -2154 4368 -2138 4402
rect -1962 4368 -1946 4402
rect -2200 4343 -2188 4359
rect -2250 4309 -2222 4320
rect -2250 4293 -2188 4309
rect -2250 4290 -2190 4293
rect -2154 4250 -2138 4284
rect -1962 4250 -1946 4284
rect -2324 4180 -2290 4232
rect -1872 4180 -1838 4232
rect -1044 4600 -948 4634
rect -654 4600 -558 4634
rect -1044 4538 -1010 4600
rect -592 4538 -558 4600
rect -970 4477 -910 4490
rect -874 4486 -858 4520
rect -682 4486 -666 4520
rect -970 4461 -908 4477
rect -970 4460 -942 4461
rect -970 4320 -960 4460
rect -920 4411 -908 4427
rect -920 4359 -910 4411
rect -874 4368 -858 4402
rect -682 4368 -666 4402
rect -920 4343 -908 4359
rect -970 4309 -942 4320
rect -970 4293 -908 4309
rect -970 4290 -910 4293
rect -874 4250 -858 4284
rect -682 4250 -666 4284
rect -1044 4180 -1010 4232
rect -592 4180 -558 4232
rect 256 4600 352 4634
rect 646 4600 742 4634
rect 256 4538 290 4600
rect 708 4538 742 4600
rect 330 4477 390 4490
rect 426 4486 442 4520
rect 618 4486 634 4520
rect 330 4461 392 4477
rect 330 4460 358 4461
rect 330 4320 340 4460
rect 380 4411 392 4427
rect 380 4359 390 4411
rect 426 4368 442 4402
rect 618 4368 634 4402
rect 380 4343 392 4359
rect 330 4309 358 4320
rect 330 4293 392 4309
rect 330 4290 390 4293
rect 426 4250 442 4284
rect 618 4250 634 4284
rect 256 4180 290 4232
rect 708 4180 742 4232
rect 1536 4600 1632 4634
rect 1926 4600 2022 4634
rect 1536 4538 1570 4600
rect 1988 4538 2022 4600
rect 1610 4477 1670 4490
rect 1706 4486 1722 4520
rect 1898 4486 1914 4520
rect 1610 4461 1672 4477
rect 1610 4460 1638 4461
rect 1610 4320 1620 4460
rect 1660 4411 1672 4427
rect 1660 4359 1670 4411
rect 1706 4368 1722 4402
rect 1898 4368 1914 4402
rect 1660 4343 1672 4359
rect 1610 4309 1638 4320
rect 1610 4293 1672 4309
rect 1610 4290 1670 4293
rect 1706 4250 1722 4284
rect 1898 4250 1914 4284
rect 1536 4180 1570 4232
rect 1988 4180 2022 4232
rect 2836 4600 2932 4634
rect 3226 4600 3322 4634
rect 2836 4538 2870 4600
rect 3288 4538 3322 4600
rect 2910 4477 2970 4490
rect 3006 4486 3022 4520
rect 3198 4486 3214 4520
rect 2910 4461 2972 4477
rect 2910 4460 2938 4461
rect 2910 4320 2920 4460
rect 2960 4411 2972 4427
rect 2960 4359 2970 4411
rect 3006 4368 3022 4402
rect 3198 4368 3214 4402
rect 2960 4343 2972 4359
rect 2910 4309 2938 4320
rect 2910 4293 2972 4309
rect 2910 4290 2970 4293
rect 3006 4250 3022 4284
rect 3198 4250 3214 4284
rect 2836 4180 2870 4232
rect 3288 4180 3322 4232
rect 4116 4600 4212 4634
rect 4506 4600 4602 4634
rect 4116 4538 4150 4600
rect 4568 4538 4602 4600
rect 4190 4477 4250 4490
rect 4286 4486 4302 4520
rect 4478 4486 4494 4520
rect 4190 4461 4252 4477
rect 4190 4460 4218 4461
rect 4190 4320 4200 4460
rect 4240 4411 4252 4427
rect 4240 4359 4250 4411
rect 4286 4368 4302 4402
rect 4478 4368 4494 4402
rect 4240 4343 4252 4359
rect 4190 4309 4218 4320
rect 4190 4293 4252 4309
rect 4190 4290 4250 4293
rect 4286 4250 4302 4284
rect 4478 4250 4494 4284
rect 4116 4180 4150 4232
rect 4568 4180 4602 4232
rect 5416 4600 5512 4634
rect 5806 4600 5902 4634
rect 5416 4538 5450 4600
rect 5868 4538 5902 4600
rect 5490 4477 5550 4490
rect 5586 4486 5602 4520
rect 5778 4486 5794 4520
rect 5490 4461 5552 4477
rect 5490 4460 5518 4461
rect 5490 4320 5500 4460
rect 5540 4411 5552 4427
rect 5540 4359 5550 4411
rect 5586 4368 5602 4402
rect 5778 4368 5794 4402
rect 5540 4343 5552 4359
rect 5490 4309 5518 4320
rect 5490 4293 5552 4309
rect 5490 4290 5550 4293
rect 5586 4250 5602 4284
rect 5778 4250 5794 4284
rect 5416 4180 5450 4232
rect 5868 4180 5902 4232
rect 6696 4600 6792 4634
rect 7086 4600 7182 4634
rect 6696 4538 6730 4600
rect 7148 4538 7182 4600
rect 6770 4477 6830 4490
rect 6866 4486 6882 4520
rect 7058 4486 7074 4520
rect 6770 4461 6832 4477
rect 6770 4460 6798 4461
rect 6770 4320 6780 4460
rect 6820 4411 6832 4427
rect 6820 4359 6830 4411
rect 6866 4368 6882 4402
rect 7058 4368 7074 4402
rect 6820 4343 6832 4359
rect 6770 4309 6798 4320
rect 6770 4293 6832 4309
rect 6770 4290 6830 4293
rect 6866 4250 6882 4284
rect 7058 4250 7074 4284
rect 6696 4180 6730 4232
rect 7148 4180 7182 4232
rect 7996 4600 8092 4634
rect 8386 4600 8482 4634
rect 7996 4538 8030 4600
rect 8448 4538 8482 4600
rect 8070 4477 8130 4490
rect 8166 4486 8182 4520
rect 8358 4486 8374 4520
rect 8070 4461 8132 4477
rect 8070 4460 8098 4461
rect 8070 4320 8080 4460
rect 8120 4411 8132 4427
rect 8120 4359 8130 4411
rect 8166 4368 8182 4402
rect 8358 4368 8374 4402
rect 8120 4343 8132 4359
rect 8070 4309 8098 4320
rect 8070 4293 8132 4309
rect 8070 4290 8130 4293
rect 8166 4250 8182 4284
rect 8358 4250 8374 4284
rect 7996 4180 8030 4232
rect 8448 4180 8482 4232
rect 9276 4600 9372 4634
rect 9666 4600 9762 4634
rect 9276 4538 9310 4600
rect 9728 4538 9762 4600
rect 9350 4477 9410 4490
rect 9446 4486 9462 4520
rect 9638 4486 9654 4520
rect 9350 4461 9412 4477
rect 9350 4460 9378 4461
rect 9350 4320 9360 4460
rect 9400 4411 9412 4427
rect 9400 4359 9410 4411
rect 9446 4368 9462 4402
rect 9638 4368 9654 4402
rect 9400 4343 9412 4359
rect 9350 4309 9378 4320
rect 9350 4293 9412 4309
rect 9350 4290 9410 4293
rect 9446 4250 9462 4284
rect 9638 4250 9654 4284
rect 9276 4180 9310 4232
rect 9728 4180 9762 4232
rect -4980 4170 9800 4180
rect -4980 4136 -4808 4170
rect -4514 4136 -3528 4170
rect -3234 4136 -2228 4170
rect -1934 4136 -948 4170
rect -654 4136 352 4170
rect 646 4136 1632 4170
rect 1926 4136 2932 4170
rect 3226 4136 4212 4170
rect 4506 4136 5512 4170
rect 5806 4136 6792 4170
rect 7086 4136 8092 4170
rect 8386 4136 9372 4170
rect 9666 4136 9800 4170
rect -4980 4100 9800 4136
rect -4980 365 -4800 4100
rect -170 2840 -70 2850
rect -170 2800 -160 2840
rect -80 2830 -70 2840
rect -80 2800 100 2830
rect -170 2790 100 2800
rect 220 2520 360 4100
rect 3430 2600 3810 2710
rect 8930 2620 9090 2710
rect 480 2560 720 2570
rect 480 2520 600 2560
rect 710 2520 720 2560
rect 480 2510 720 2520
rect -4385 1800 -3950 1820
rect -4400 1750 -3950 1800
rect -4400 1500 -4350 1750
rect -4200 1710 -3950 1750
rect -4200 1500 -4150 1710
rect -4400 1450 -4150 1500
rect -5065 -2385 -4755 55
rect -4385 90 -4175 1450
rect -4020 1300 -3940 1320
rect -4020 1240 -4000 1300
rect -3960 1240 -3940 1300
rect -4020 1220 -3940 1240
rect -3000 1300 -2900 1320
rect -3000 1240 -2980 1300
rect -2920 1240 -2900 1300
rect -3000 1220 -2900 1240
rect -1940 1300 -1840 1320
rect -1940 1240 -1920 1300
rect -1860 1240 -1840 1300
rect -1940 1220 -1840 1240
rect -920 1300 -820 1320
rect -920 1240 -900 1300
rect -840 1240 -820 1300
rect -920 1220 -820 1240
rect -4065 549 -3755 715
rect 90 680 385 790
rect 90 660 200 680
rect -4065 251 -4059 549
rect -3761 251 -3755 549
rect -4065 245 -3755 251
rect 3440 90 3610 2600
rect 5820 2130 5830 2190
rect 8210 90 8390 580
rect -4385 -90 8400 90
rect -4385 -120 -3780 -90
rect -450 -150 850 -90
rect 4250 -160 4870 -90
rect 110 -1760 380 -1750
rect 110 -1800 120 -1760
rect 180 -1790 380 -1760
rect 180 -1800 190 -1790
rect 110 -1810 190 -1800
rect 260 -2350 350 -1860
rect -5065 -2450 -3680 -2385
rect -650 -2450 1350 -2350
rect 4110 -2450 4940 -2400
rect 8570 -2450 8680 1630
rect 8930 1570 9070 1650
rect -5065 -2540 8700 -2450
rect -5065 -2660 9420 -2540
rect -5065 -2670 8700 -2660
rect -5065 -2695 -3680 -2670
rect -3990 -5600 -3680 -2695
rect 7220 -4210 7320 -3220
rect 7210 -4290 7320 -4210
rect 7380 -3890 7500 -2670
rect 8570 -2680 8680 -2670
rect 11160 -3360 12140 -3300
rect 7380 -4350 7480 -3890
rect 11160 -4090 11220 -3360
rect 12410 -3390 12490 -3290
rect 12400 -3820 12480 -3800
rect 12400 -3900 12420 -3820
rect 12460 -3900 12480 -3820
rect 12400 -3920 12480 -3900
rect 11100 -4096 11280 -4090
rect 8100 -4310 8190 -4210
rect 11100 -4264 11106 -4096
rect 11274 -4264 11280 -4096
rect 7380 -4600 7500 -4350
rect 8100 -4590 8200 -4310
rect 11100 -4590 11280 -4264
rect 11540 -4206 11980 -4200
rect 11540 -4314 11566 -4206
rect 11674 -4314 11980 -4206
rect 11540 -4400 11980 -4314
rect 12410 -4430 12490 -4350
rect 7920 -4690 8200 -4590
rect 10230 -4800 16130 -4590
rect 12070 -4880 12550 -4800
rect 7320 -4940 7410 -4930
rect 5980 -5600 6120 -5550
rect -4000 -5680 -3680 -5600
rect -4000 -5800 4200 -5680
rect 4460 -5700 7680 -5600
rect 4840 -5780 4900 -5700
rect 5340 -5780 5400 -5700
rect 5860 -5780 5920 -5700
rect 6380 -5780 6440 -5700
rect 6900 -5780 6960 -5700
rect 7420 -5780 7480 -5700
rect -4000 -5880 -3680 -5800
rect 7560 -5840 7680 -5700
rect -4000 -7120 -3690 -5880
rect 7560 -5920 8200 -5840
rect 7560 -6100 7800 -5920
rect 7560 -6180 7780 -6100
rect 4580 -7120 4640 -6980
rect 5100 -7120 5160 -6960
rect 5600 -7120 5660 -6960
rect 6120 -7120 6180 -6960
rect 6640 -7120 6700 -6940
rect 7160 -7120 7220 -6940
rect 7640 -7120 7780 -6860
rect 8640 -7100 8740 -7080
rect 8640 -7120 9890 -7100
rect -4000 -7150 9890 -7120
rect 11560 -7150 12760 -7070
rect -4000 -7240 15540 -7150
rect -4000 -7300 8640 -7240
rect 9780 -7310 15540 -7240
rect 11600 -7381 11750 -7310
rect 11600 -7519 11606 -7381
rect 11744 -7519 11750 -7381
rect 11600 -7525 11750 -7519
rect 9000 -7580 9100 -7570
rect 8840 -7620 9020 -7580
rect 9080 -7620 9100 -7580
rect 9000 -7630 9100 -7620
rect 9400 -7580 9670 -7570
rect 9400 -7620 9610 -7580
rect 9650 -7620 9670 -7580
rect 9400 -7630 9670 -7620
<< viali >>
rect -4350 5130 -4310 5180
rect -4820 4960 -4780 5100
rect -4340 4880 -4300 4930
rect -3428 5126 -3252 5160
rect -3530 5067 -3512 5100
rect -3512 5067 -3490 5100
rect -3530 4983 -3490 5067
rect -3428 5008 -3252 5042
rect -3530 4960 -3512 4983
rect -3512 4960 -3490 4983
rect -3428 4890 -3252 4924
rect -3060 5130 -3020 5180
rect -3050 4880 -3010 4930
rect -2138 5126 -1962 5160
rect -2240 5067 -2222 5100
rect -2222 5067 -2200 5100
rect -2240 4983 -2200 5067
rect -2138 5008 -1962 5042
rect -2240 4960 -2222 4983
rect -2222 4960 -2200 4983
rect -2138 4890 -1962 4924
rect -1770 5130 -1730 5180
rect -1760 4880 -1720 4930
rect -848 5126 -672 5160
rect -950 5067 -932 5100
rect -932 5067 -910 5100
rect -950 4983 -910 5067
rect -848 5008 -672 5042
rect -950 4960 -932 4983
rect -932 4960 -910 4983
rect -848 4890 -672 4924
rect -480 5130 -440 5180
rect -470 4880 -430 4930
rect 442 5126 618 5160
rect 340 5067 358 5100
rect 358 5067 380 5100
rect 340 4983 380 5067
rect 442 5008 618 5042
rect 340 4960 358 4983
rect 358 4960 380 4983
rect 442 4890 618 4924
rect 810 5130 850 5180
rect 820 4880 860 4930
rect 1732 5126 1908 5160
rect 1630 5067 1648 5100
rect 1648 5067 1670 5100
rect 1630 4983 1670 5067
rect 1732 5008 1908 5042
rect 1630 4960 1648 4983
rect 1648 4960 1670 4983
rect 1732 4890 1908 4924
rect 2100 5130 2140 5180
rect 2110 4880 2150 4930
rect 3022 5126 3198 5160
rect 2920 5067 2938 5100
rect 2938 5067 2960 5100
rect 2920 4983 2960 5067
rect 3022 5008 3198 5042
rect 2920 4960 2938 4983
rect 2938 4960 2960 4983
rect 3022 4890 3198 4924
rect 3390 5130 3430 5180
rect 3400 4880 3440 4930
rect 4312 5126 4488 5160
rect 4210 5067 4228 5100
rect 4228 5067 4250 5100
rect 4210 4983 4250 5067
rect 4312 5008 4488 5042
rect 4210 4960 4228 4983
rect 4228 4960 4250 4983
rect 4312 4890 4488 4924
rect 4680 5130 4720 5180
rect 4690 4880 4730 4930
rect 5602 5126 5778 5160
rect 5500 5067 5518 5100
rect 5518 5067 5540 5100
rect 5500 4983 5540 5067
rect 5602 5008 5778 5042
rect 5500 4960 5518 4983
rect 5518 4960 5540 4983
rect 5602 4890 5778 4924
rect 5970 5130 6010 5180
rect 5980 4880 6020 4930
rect 6892 5126 7068 5160
rect 6790 5067 6808 5100
rect 6808 5067 6830 5100
rect 6790 4983 6830 5067
rect 6892 5008 7068 5042
rect 6790 4960 6808 4983
rect 6808 4960 6830 4983
rect 6892 4890 7068 4924
rect 7260 5130 7300 5180
rect 7270 4880 7310 4930
rect 8182 5126 8358 5160
rect 8080 5067 8098 5100
rect 8098 5067 8120 5100
rect 8080 4983 8120 5067
rect 8182 5008 8358 5042
rect 8080 4960 8098 4983
rect 8098 4960 8120 4983
rect 8182 4890 8358 4924
rect 8550 5130 8590 5180
rect 8560 4880 8600 4930
rect 9472 5126 9648 5160
rect 9370 5067 9388 5100
rect 9388 5067 9410 5100
rect 9370 4983 9410 5067
rect 9472 5008 9648 5042
rect 9370 4960 9388 4983
rect 9388 4960 9410 4983
rect 9472 4890 9648 4924
rect 9840 5130 9880 5180
rect 9850 4880 9890 4930
rect -4718 4486 -4542 4520
rect -4820 4427 -4802 4460
rect -4802 4427 -4780 4460
rect -4820 4343 -4780 4427
rect -4718 4368 -4542 4402
rect -4820 4320 -4802 4343
rect -4802 4320 -4780 4343
rect -4718 4250 -4542 4284
rect -3438 4486 -3262 4520
rect -3540 4427 -3522 4460
rect -3522 4427 -3500 4460
rect -3540 4343 -3500 4427
rect -3438 4368 -3262 4402
rect -3540 4320 -3522 4343
rect -3522 4320 -3500 4343
rect -3438 4250 -3262 4284
rect -2138 4486 -1962 4520
rect -2240 4427 -2222 4460
rect -2222 4427 -2200 4460
rect -2240 4343 -2200 4427
rect -2138 4368 -1962 4402
rect -2240 4320 -2222 4343
rect -2222 4320 -2200 4343
rect -2138 4250 -1962 4284
rect -858 4486 -682 4520
rect -960 4427 -942 4460
rect -942 4427 -920 4460
rect -960 4343 -920 4427
rect -858 4368 -682 4402
rect -960 4320 -942 4343
rect -942 4320 -920 4343
rect -858 4250 -682 4284
rect 442 4486 618 4520
rect 340 4427 358 4460
rect 358 4427 380 4460
rect 340 4343 380 4427
rect 442 4368 618 4402
rect 340 4320 358 4343
rect 358 4320 380 4343
rect 442 4250 618 4284
rect 1722 4486 1898 4520
rect 1620 4427 1638 4460
rect 1638 4427 1660 4460
rect 1620 4343 1660 4427
rect 1722 4368 1898 4402
rect 1620 4320 1638 4343
rect 1638 4320 1660 4343
rect 1722 4250 1898 4284
rect 3022 4486 3198 4520
rect 2920 4427 2938 4460
rect 2938 4427 2960 4460
rect 2920 4343 2960 4427
rect 3022 4368 3198 4402
rect 2920 4320 2938 4343
rect 2938 4320 2960 4343
rect 3022 4250 3198 4284
rect 4302 4486 4478 4520
rect 4200 4427 4218 4460
rect 4218 4427 4240 4460
rect 4200 4343 4240 4427
rect 4302 4368 4478 4402
rect 4200 4320 4218 4343
rect 4218 4320 4240 4343
rect 4302 4250 4478 4284
rect 5602 4486 5778 4520
rect 5500 4427 5518 4460
rect 5518 4427 5540 4460
rect 5500 4343 5540 4427
rect 5602 4368 5778 4402
rect 5500 4320 5518 4343
rect 5518 4320 5540 4343
rect 5602 4250 5778 4284
rect 6882 4486 7058 4520
rect 6780 4427 6798 4460
rect 6798 4427 6820 4460
rect 6780 4343 6820 4427
rect 6882 4368 7058 4402
rect 6780 4320 6798 4343
rect 6798 4320 6820 4343
rect 6882 4250 7058 4284
rect 8182 4486 8358 4520
rect 8080 4427 8098 4460
rect 8098 4427 8120 4460
rect 8080 4343 8120 4427
rect 8182 4368 8358 4402
rect 8080 4320 8098 4343
rect 8098 4320 8120 4343
rect 8182 4250 8358 4284
rect 9462 4486 9638 4520
rect 9360 4427 9378 4460
rect 9378 4427 9400 4460
rect 9360 4343 9400 4427
rect 9462 4368 9638 4402
rect 9360 4320 9378 4343
rect 9378 4320 9400 4343
rect 9462 4250 9638 4284
rect -160 2800 -80 2840
rect 600 2520 710 2560
rect -4350 1500 -4200 1750
rect -5065 55 -4755 365
rect -4000 1240 -3960 1300
rect -2980 1240 -2920 1300
rect -1920 1240 -1860 1300
rect -900 1240 -840 1300
rect 385 680 495 790
rect -4059 251 -3761 549
rect 3720 2130 3780 2190
rect 4770 2130 4830 2190
rect 5830 2130 5890 2190
rect 6860 2130 6920 2190
rect 7910 2130 7970 2190
rect 8210 580 8390 760
rect 120 -1800 180 -1760
rect 9420 -2660 9540 -2540
rect 7220 -3220 7320 -3120
rect 12420 -3900 12460 -3820
rect 13500 -3870 13560 -3810
rect 8190 -4310 8290 -4210
rect 11106 -4264 11274 -4096
rect 11566 -4314 11674 -4206
rect 7320 -4930 7420 -4830
rect 5980 -5550 6120 -5410
rect 11606 -7519 11744 -7381
rect 9020 -7620 9080 -7580
rect 9610 -7620 9650 -7580
<< metal1 >>
rect -7690 7450 9390 7510
rect -7810 6890 -7750 6896
rect -7690 6890 -7630 7450
rect -7750 6830 -7630 6890
rect -7570 7350 9110 7410
rect -7810 6824 -7750 6830
rect -7690 6770 -7630 6776
rect -7570 6770 -7510 7350
rect -7630 6710 -7510 6770
rect -7470 7250 8090 7310
rect -7690 6704 -7630 6710
rect -7470 6650 -7410 7250
rect -7576 6590 -7570 6650
rect -7510 6590 -7410 6650
rect -7330 7150 7770 7210
rect -7330 6550 -7270 7150
rect -7476 6490 -7470 6550
rect -7410 6490 -7270 6550
rect -7210 7050 6810 7110
rect -7210 6450 -7150 7050
rect -7356 6390 -7350 6450
rect -7290 6390 -7150 6450
rect -7090 6950 6510 7010
rect -7090 6350 -7030 6950
rect -7236 6290 -7230 6350
rect -7170 6290 -7030 6350
rect -6990 6850 5510 6910
rect -6990 6250 -6930 6850
rect -7096 6190 -7090 6250
rect -7030 6190 -6930 6250
rect -6870 6750 5210 6810
rect -6870 6150 -6810 6750
rect -6976 6090 -6970 6150
rect -6910 6090 -6810 6150
rect -6750 6650 3950 6710
rect -6750 6050 -6690 6650
rect -6856 5990 -6850 6050
rect -6790 5990 -6690 6050
rect -6630 6550 2930 6610
rect -6630 5950 -6570 6550
rect -6736 5890 -6730 5950
rect -6670 5890 -6570 5950
rect -6510 6450 2630 6510
rect -6510 5850 -6450 6450
rect -6596 5790 -6590 5850
rect -6530 5790 -6450 5850
rect -6410 6330 1650 6390
rect -6476 5690 -6470 5750
rect -6410 5690 -6350 6330
rect -6290 6210 1350 6270
rect -6356 5590 -6350 5650
rect -6290 5590 -6230 6210
rect -6190 6110 370 6170
rect -6190 5516 -6130 6110
rect -6250 5510 -6130 5516
rect -6190 5450 -6130 5510
rect -6070 6010 70 6070
rect -6250 5444 -6190 5450
rect -6136 5330 -6130 5390
rect -6070 5330 -6010 6010
rect -5950 5890 -930 5950
rect -6016 5230 -6010 5290
rect -5950 5230 -5890 5890
rect -5850 5770 -1230 5830
rect -5916 5130 -5910 5190
rect -5850 5130 -5790 5770
rect -5750 5650 -2210 5710
rect -5750 5090 -5690 5650
rect -5796 5030 -5790 5090
rect -5730 5030 -5690 5090
rect -5630 5530 -2550 5590
rect -5696 4910 -5690 4970
rect -5630 4910 -5570 5530
rect -5510 5430 -3490 5490
rect -5510 4870 -5450 5430
rect -5596 4810 -5590 4870
rect -5530 4810 -5450 4870
rect -5390 5310 -3830 5370
rect -5390 4770 -5330 5310
rect -4486 5181 -4434 5187
rect -4630 5130 -4486 5180
rect -4830 5100 -4770 5130
rect -4360 5180 -4300 5200
rect -4434 5130 -4350 5180
rect -4310 5130 -4300 5180
rect -4486 5123 -4434 5129
rect -4360 5110 -4300 5130
rect -5250 5050 -5190 5056
rect -4830 5050 -4820 5100
rect -5190 4990 -4820 5050
rect -5250 4984 -5190 4990
rect -4830 4960 -4820 4990
rect -4780 4960 -4770 5100
rect -4630 5000 -4020 5050
rect -4830 4930 -4770 4960
rect -4350 4930 -4290 4950
rect -4630 4880 -4340 4930
rect -4300 4880 -4290 4930
rect -5476 4710 -5470 4770
rect -5410 4710 -5330 4770
rect -4465 4540 -4415 4880
rect -4350 4860 -4290 4880
rect -4610 4526 -4150 4540
rect -4730 4520 -4150 4526
rect -4830 4460 -4770 4490
rect -4730 4486 -4718 4520
rect -4542 4490 -4150 4520
rect -4542 4486 -4530 4490
rect -4730 4480 -4530 4486
rect -4830 4410 -4820 4460
rect -5250 4350 -4820 4410
rect -5250 3890 -5190 4350
rect -4830 4320 -4820 4350
rect -4780 4320 -4770 4460
rect -4310 4411 -4240 4420
rect -4310 4410 -4301 4411
rect -4620 4408 -4301 4410
rect -4730 4402 -4301 4408
rect -4730 4368 -4718 4402
rect -4542 4368 -4301 4402
rect -4730 4362 -4301 4368
rect -4620 4360 -4301 4362
rect -4310 4359 -4301 4360
rect -4249 4359 -4240 4411
rect -4310 4350 -4240 4359
rect -4830 4290 -4770 4320
rect -4730 4284 -4530 4290
rect -4730 4250 -4718 4284
rect -4542 4280 -4530 4284
rect -4200 4280 -4150 4490
rect -4542 4250 -4150 4280
rect -4730 4244 -4150 4250
rect -4620 4230 -4150 4244
rect -4070 4100 -4020 5000
rect -3890 4390 -3830 5310
rect -3550 5130 -3490 5430
rect -3210 5306 -3158 5312
rect -3210 5248 -3158 5254
rect -3209 5180 -3159 5248
rect -3070 5180 -3010 5200
rect -3340 5166 -3060 5180
rect -3440 5160 -3060 5166
rect -3550 5100 -3480 5130
rect -3440 5126 -3428 5160
rect -3252 5130 -3060 5160
rect -3020 5130 -3010 5180
rect -3252 5126 -3240 5130
rect -3440 5120 -3240 5126
rect -3070 5110 -3010 5130
rect -3550 4960 -3530 5100
rect -3490 4960 -3480 5100
rect -3340 5048 -2730 5050
rect -3440 5042 -2730 5048
rect -3440 5008 -3428 5042
rect -3252 5008 -2730 5042
rect -3440 5002 -2730 5008
rect -3340 5000 -2730 5002
rect -3550 4930 -3480 4960
rect -3060 4930 -3000 4950
rect -3440 4924 -3050 4930
rect -3440 4890 -3428 4924
rect -3252 4890 -3050 4924
rect -3440 4884 -3050 4890
rect -3340 4880 -3050 4884
rect -3010 4880 -3000 4930
rect -3225 4540 -3175 4880
rect -3060 4860 -3000 4880
rect -3330 4526 -2870 4540
rect -3450 4520 -2870 4526
rect -3550 4460 -3490 4490
rect -3450 4486 -3438 4520
rect -3262 4490 -2870 4520
rect -3262 4486 -3250 4490
rect -3450 4480 -3250 4486
rect -3550 4390 -3540 4460
rect -3890 4330 -3540 4390
rect -3550 4320 -3540 4330
rect -3500 4320 -3490 4460
rect -3030 4411 -2960 4420
rect -3030 4410 -3021 4411
rect -3340 4408 -3021 4410
rect -3450 4402 -3021 4408
rect -3450 4368 -3438 4402
rect -3262 4368 -3021 4402
rect -3450 4362 -3021 4368
rect -3340 4360 -3021 4362
rect -3030 4359 -3021 4360
rect -2969 4359 -2960 4411
rect -3030 4350 -2960 4359
rect -3550 4290 -3490 4320
rect -3450 4284 -3250 4290
rect -3450 4250 -3438 4284
rect -3262 4280 -3250 4284
rect -2920 4280 -2870 4490
rect -3262 4250 -2870 4280
rect -3450 4244 -2870 4250
rect -3340 4230 -2870 4244
rect -2780 4100 -2730 5000
rect -2610 4410 -2550 5530
rect -2270 5130 -2210 5650
rect -1930 5482 -1878 5488
rect -1930 5424 -1878 5430
rect -1929 5180 -1879 5424
rect -1780 5180 -1720 5200
rect -2050 5166 -1770 5180
rect -2150 5160 -1770 5166
rect -2270 5100 -2190 5130
rect -2150 5126 -2138 5160
rect -1962 5130 -1770 5160
rect -1730 5130 -1720 5180
rect -1962 5126 -1950 5130
rect -2150 5120 -1950 5126
rect -1780 5110 -1720 5130
rect -2270 4960 -2240 5100
rect -2200 4960 -2190 5100
rect -2050 5048 -1440 5050
rect -2150 5042 -1440 5048
rect -2150 5008 -2138 5042
rect -1962 5008 -1440 5042
rect -2150 5002 -1440 5008
rect -2050 5000 -1440 5002
rect -2270 4950 -2190 4960
rect -2250 4930 -2190 4950
rect -1770 4930 -1710 4950
rect -2150 4924 -1760 4930
rect -2150 4890 -2138 4924
rect -1962 4890 -1760 4924
rect -2150 4884 -1760 4890
rect -2050 4880 -1760 4884
rect -1720 4880 -1710 4930
rect -1936 4540 -1872 4880
rect -1770 4860 -1710 4880
rect -2030 4526 -1570 4540
rect -2150 4520 -1570 4526
rect -2250 4460 -2190 4490
rect -2150 4486 -2138 4520
rect -1962 4490 -1570 4520
rect -1962 4486 -1950 4490
rect -2150 4480 -1950 4486
rect -2250 4410 -2240 4460
rect -2610 4350 -2240 4410
rect -2250 4320 -2240 4350
rect -2200 4320 -2190 4460
rect -1730 4411 -1660 4420
rect -1730 4410 -1721 4411
rect -2040 4408 -1721 4410
rect -2150 4402 -1721 4408
rect -2150 4368 -2138 4402
rect -1962 4368 -1721 4402
rect -2150 4362 -1721 4368
rect -2040 4360 -1721 4362
rect -1730 4359 -1721 4360
rect -1669 4359 -1660 4411
rect -1730 4350 -1660 4359
rect -2250 4290 -2190 4320
rect -2150 4284 -1950 4290
rect -2150 4250 -2138 4284
rect -1962 4280 -1950 4284
rect -1620 4280 -1570 4490
rect -1962 4250 -1570 4280
rect -2150 4244 -1570 4250
rect -2040 4230 -1570 4244
rect -1490 4100 -1440 5000
rect -1290 4410 -1230 5770
rect -990 5130 -930 5890
rect -650 5594 -598 5600
rect -650 5536 -598 5542
rect -649 5180 -599 5536
rect -490 5180 -430 5200
rect -760 5166 -480 5180
rect -860 5160 -480 5166
rect -990 5100 -900 5130
rect -860 5126 -848 5160
rect -672 5130 -480 5160
rect -440 5130 -430 5180
rect -672 5126 -660 5130
rect -860 5120 -660 5126
rect -490 5110 -430 5130
rect -990 4960 -950 5100
rect -910 4960 -900 5100
rect -760 5048 -150 5050
rect -860 5042 -150 5048
rect -860 5008 -848 5042
rect -672 5008 -150 5042
rect -860 5002 -150 5008
rect -760 5000 -150 5002
rect -990 4930 -900 4960
rect -480 4930 -420 4950
rect -860 4924 -470 4930
rect -860 4890 -848 4924
rect -672 4890 -470 4924
rect -860 4884 -470 4890
rect -760 4880 -470 4884
rect -430 4880 -420 4930
rect -640 4540 -576 4880
rect -480 4860 -420 4880
rect -750 4526 -290 4540
rect -870 4520 -290 4526
rect -970 4460 -910 4490
rect -870 4486 -858 4520
rect -682 4490 -290 4520
rect -682 4486 -670 4490
rect -870 4480 -670 4486
rect -970 4410 -960 4460
rect -1290 4350 -960 4410
rect -970 4320 -960 4350
rect -920 4320 -910 4460
rect -450 4411 -380 4420
rect -450 4410 -441 4411
rect -760 4408 -441 4410
rect -870 4402 -441 4408
rect -870 4368 -858 4402
rect -682 4368 -441 4402
rect -870 4362 -441 4368
rect -760 4360 -441 4362
rect -450 4359 -441 4360
rect -389 4359 -380 4411
rect -450 4350 -380 4359
rect -970 4290 -910 4320
rect -870 4284 -670 4290
rect -870 4250 -858 4284
rect -682 4280 -670 4284
rect -340 4280 -290 4490
rect -682 4250 -290 4280
rect -870 4244 -290 4250
rect -760 4230 -290 4244
rect -200 4100 -150 5000
rect 10 4430 70 6010
rect 310 5130 370 6110
rect 640 5350 646 5402
rect 698 5350 704 5402
rect 647 5180 697 5350
rect 800 5180 860 5200
rect 530 5166 810 5180
rect 430 5160 810 5166
rect 310 5100 390 5130
rect 430 5126 442 5160
rect 618 5130 810 5160
rect 850 5130 860 5180
rect 618 5126 630 5130
rect 430 5120 630 5126
rect 800 5110 860 5130
rect 310 4960 340 5100
rect 380 4960 390 5100
rect 530 5048 1140 5050
rect 430 5042 1140 5048
rect 430 5008 442 5042
rect 618 5008 1140 5042
rect 430 5002 1140 5008
rect 530 5000 1140 5002
rect 310 4930 390 4960
rect 810 4930 870 4950
rect 430 4924 820 4930
rect 430 4890 442 4924
rect 618 4890 820 4924
rect 430 4884 820 4890
rect 530 4880 820 4884
rect 860 4880 870 4930
rect 688 4540 752 4880
rect 810 4860 870 4880
rect 550 4526 1010 4540
rect 430 4520 1010 4526
rect 330 4460 390 4490
rect 430 4486 442 4520
rect 618 4490 1010 4520
rect 618 4486 630 4490
rect 430 4480 630 4486
rect 330 4430 340 4460
rect 10 4370 340 4430
rect 330 4320 340 4370
rect 380 4320 390 4460
rect 850 4411 920 4420
rect 850 4410 859 4411
rect 540 4408 859 4410
rect 430 4402 859 4408
rect 430 4368 442 4402
rect 618 4368 859 4402
rect 430 4362 859 4368
rect 540 4360 859 4362
rect 850 4359 859 4360
rect 911 4359 920 4411
rect 850 4350 920 4359
rect 330 4290 390 4320
rect 430 4284 630 4290
rect 430 4250 442 4284
rect 618 4280 630 4284
rect 960 4280 1010 4490
rect 618 4250 1010 4280
rect 430 4244 1010 4250
rect 540 4230 1010 4244
rect 1090 4100 1140 5000
rect 1290 4410 1350 6210
rect 1590 5130 1650 6330
rect 1926 5562 1978 5568
rect 1926 5504 1978 5510
rect 1927 5180 1977 5504
rect 2090 5180 2150 5200
rect 1820 5166 2100 5180
rect 1720 5160 2100 5166
rect 1590 5100 1680 5130
rect 1720 5126 1732 5160
rect 1908 5130 2100 5160
rect 2140 5130 2150 5180
rect 1908 5126 1920 5130
rect 1720 5120 1920 5126
rect 2090 5110 2150 5130
rect 1590 4960 1630 5100
rect 1670 4960 1680 5100
rect 1820 5048 2430 5050
rect 1720 5042 2430 5048
rect 1720 5008 1732 5042
rect 1908 5008 2430 5042
rect 1720 5002 2430 5008
rect 1820 5000 2430 5002
rect 1590 4930 1680 4960
rect 2100 4930 2160 4950
rect 1720 4924 2110 4930
rect 1720 4890 1732 4924
rect 1908 4890 2110 4924
rect 1720 4884 2110 4890
rect 1820 4880 2110 4884
rect 2150 4880 2160 4930
rect 1984 4540 2048 4880
rect 2100 4860 2160 4880
rect 1830 4526 2290 4540
rect 1710 4520 2290 4526
rect 1610 4460 1670 4490
rect 1710 4486 1722 4520
rect 1898 4490 2290 4520
rect 1898 4486 1910 4490
rect 1710 4480 1910 4486
rect 1610 4410 1620 4460
rect 1290 4350 1620 4410
rect 1610 4320 1620 4350
rect 1660 4320 1670 4460
rect 2130 4411 2200 4420
rect 2130 4410 2139 4411
rect 1820 4408 2139 4410
rect 1710 4402 2139 4408
rect 1710 4368 1722 4402
rect 1898 4368 2139 4402
rect 1710 4362 2139 4368
rect 1820 4360 2139 4362
rect 2130 4359 2139 4360
rect 2191 4359 2200 4411
rect 2130 4350 2200 4359
rect 1610 4290 1670 4320
rect 1710 4284 1910 4290
rect 1710 4250 1722 4284
rect 1898 4280 1910 4284
rect 2240 4280 2290 4490
rect 1898 4250 2290 4280
rect 1710 4244 2290 4250
rect 1820 4230 2290 4244
rect 2380 4100 2430 5000
rect 2570 4410 2630 6450
rect 2870 5130 2930 6550
rect 3238 5738 3290 5744
rect 3238 5680 3290 5686
rect 3239 5180 3289 5680
rect 3380 5180 3440 5200
rect 3110 5166 3390 5180
rect 3010 5160 3390 5166
rect 2870 5100 2970 5130
rect 3010 5126 3022 5160
rect 3198 5130 3390 5160
rect 3430 5130 3440 5180
rect 3198 5126 3210 5130
rect 3010 5120 3210 5126
rect 3380 5110 3440 5130
rect 2870 4960 2920 5100
rect 2960 4960 2970 5100
rect 3110 5048 3720 5050
rect 3010 5042 3720 5048
rect 3010 5008 3022 5042
rect 3198 5008 3720 5042
rect 3010 5002 3720 5008
rect 3110 5000 3720 5002
rect 2870 4930 2970 4960
rect 3390 4930 3450 4950
rect 3010 4924 3400 4930
rect 3010 4890 3022 4924
rect 3198 4890 3400 4924
rect 3010 4884 3400 4890
rect 3110 4880 3400 4884
rect 3440 4880 3450 4930
rect 3264 4540 3328 4880
rect 3390 4860 3450 4880
rect 3130 4526 3590 4540
rect 3010 4520 3590 4526
rect 2910 4460 2970 4490
rect 3010 4486 3022 4520
rect 3198 4490 3590 4520
rect 3198 4486 3210 4490
rect 3010 4480 3210 4486
rect 2910 4410 2920 4460
rect 2570 4350 2920 4410
rect 2910 4320 2920 4350
rect 2960 4320 2970 4460
rect 3430 4411 3500 4420
rect 3430 4410 3439 4411
rect 3120 4408 3439 4410
rect 3010 4402 3439 4408
rect 3010 4368 3022 4402
rect 3198 4368 3439 4402
rect 3010 4362 3439 4368
rect 3120 4360 3439 4362
rect 3430 4359 3439 4360
rect 3491 4359 3500 4411
rect 3430 4350 3500 4359
rect 2910 4290 2970 4320
rect 3010 4284 3210 4290
rect 3010 4250 3022 4284
rect 3198 4280 3210 4284
rect 3540 4280 3590 4490
rect 3198 4250 3590 4280
rect 3010 4244 3590 4250
rect 3120 4230 3590 4244
rect 3670 4100 3720 5000
rect 3890 4410 3950 6650
rect 4534 5978 4586 5984
rect 4534 5920 4586 5926
rect 4170 5376 4176 5440
rect 4240 5376 4246 5440
rect 4176 5130 4240 5376
rect 4535 5180 4585 5920
rect 4670 5180 4730 5200
rect 4400 5166 4680 5180
rect 4300 5160 4680 5166
rect 4176 5100 4260 5130
rect 4300 5126 4312 5160
rect 4488 5130 4680 5160
rect 4720 5130 4730 5180
rect 4488 5126 4500 5130
rect 4300 5120 4500 5126
rect 4670 5110 4730 5130
rect 4176 4960 4210 5100
rect 4250 4960 4260 5100
rect 4400 5048 5010 5050
rect 4300 5042 5010 5048
rect 4300 5008 4312 5042
rect 4488 5008 5010 5042
rect 4300 5002 5010 5008
rect 4400 5000 5010 5002
rect 4200 4930 4260 4960
rect 4680 4930 4740 4950
rect 4300 4924 4690 4930
rect 4300 4890 4312 4924
rect 4488 4890 4690 4924
rect 4300 4884 4690 4890
rect 4400 4880 4690 4884
rect 4730 4880 4740 4930
rect 4576 4540 4640 4880
rect 4680 4860 4740 4880
rect 4410 4526 4870 4540
rect 4290 4520 4870 4526
rect 4190 4460 4250 4490
rect 4290 4486 4302 4520
rect 4478 4490 4870 4520
rect 4478 4486 4490 4490
rect 4290 4480 4490 4486
rect 4190 4410 4200 4460
rect 3890 4350 4200 4410
rect 4190 4320 4200 4350
rect 4240 4320 4250 4460
rect 4710 4411 4780 4420
rect 4710 4410 4719 4411
rect 4400 4408 4719 4410
rect 4290 4402 4719 4408
rect 4290 4368 4302 4402
rect 4478 4368 4719 4402
rect 4290 4362 4719 4368
rect 4400 4360 4719 4362
rect 4710 4359 4719 4360
rect 4771 4359 4780 4411
rect 4710 4350 4780 4359
rect 4190 4290 4250 4320
rect 4290 4284 4490 4290
rect 4290 4250 4302 4284
rect 4478 4280 4490 4284
rect 4820 4280 4870 4490
rect 4478 4250 4870 4280
rect 4290 4244 4870 4250
rect 4400 4230 4870 4244
rect 4960 4100 5010 5000
rect 5150 4410 5210 6750
rect 5450 5130 5510 6850
rect 5814 6186 5866 6192
rect 5814 6128 5866 6134
rect 5815 5180 5865 6128
rect 5960 5180 6020 5200
rect 5690 5166 5970 5180
rect 5590 5160 5970 5166
rect 5450 5100 5550 5130
rect 5590 5126 5602 5160
rect 5778 5130 5970 5160
rect 6010 5130 6020 5180
rect 5778 5126 5790 5130
rect 5590 5120 5790 5126
rect 5960 5110 6020 5130
rect 5450 4960 5500 5100
rect 5540 4960 5550 5100
rect 5690 5048 6300 5050
rect 5590 5042 6300 5048
rect 5590 5008 5602 5042
rect 5778 5008 6300 5042
rect 5590 5002 6300 5008
rect 5690 5000 6300 5002
rect 5450 4950 5550 4960
rect 5490 4930 5550 4950
rect 5970 4930 6030 4950
rect 5590 4924 5980 4930
rect 5590 4890 5602 4924
rect 5778 4890 5980 4924
rect 5590 4884 5980 4890
rect 5690 4880 5980 4884
rect 6020 4880 6030 4930
rect 5856 4540 5920 4880
rect 5970 4860 6030 4880
rect 5710 4526 6170 4540
rect 5590 4520 6170 4526
rect 5490 4460 5550 4490
rect 5590 4486 5602 4520
rect 5778 4490 6170 4520
rect 5778 4486 5790 4490
rect 5590 4480 5790 4486
rect 5490 4410 5500 4460
rect 5150 4350 5500 4410
rect 5490 4320 5500 4350
rect 5540 4320 5550 4460
rect 6010 4411 6080 4420
rect 6010 4410 6019 4411
rect 5700 4408 6019 4410
rect 5590 4402 6019 4408
rect 5590 4368 5602 4402
rect 5778 4368 6019 4402
rect 5590 4362 6019 4368
rect 5700 4360 6019 4362
rect 6010 4359 6019 4360
rect 6071 4359 6080 4411
rect 6010 4350 6080 4359
rect 5490 4290 5550 4320
rect 5590 4284 5790 4290
rect 5590 4250 5602 4284
rect 5778 4280 5790 4284
rect 6120 4280 6170 4490
rect 5778 4250 6170 4280
rect 5590 4244 6170 4250
rect 5700 4230 6170 4244
rect 6250 4100 6300 5000
rect 6450 4410 6510 6950
rect 6750 5130 6810 7050
rect 7110 5466 7162 5472
rect 7110 5408 7162 5414
rect 7111 5180 7161 5408
rect 7250 5180 7310 5200
rect 6980 5166 7260 5180
rect 6880 5160 7260 5166
rect 6750 5100 6840 5130
rect 6880 5126 6892 5160
rect 7068 5130 7260 5160
rect 7300 5130 7310 5180
rect 7068 5126 7080 5130
rect 6880 5120 7080 5126
rect 7250 5110 7310 5130
rect 6750 4960 6790 5100
rect 6830 4960 6840 5100
rect 6980 5048 7590 5050
rect 6880 5042 7590 5048
rect 6880 5008 6892 5042
rect 7068 5008 7590 5042
rect 6880 5002 7590 5008
rect 6980 5000 7590 5002
rect 6750 4930 6840 4960
rect 7260 4930 7320 4950
rect 6880 4924 7270 4930
rect 6880 4890 6892 4924
rect 7068 4890 7270 4924
rect 6880 4884 7270 4890
rect 6980 4880 7270 4884
rect 7310 4880 7320 4930
rect 7152 4540 7216 4880
rect 7260 4860 7320 4880
rect 6990 4526 7450 4540
rect 6870 4520 7450 4526
rect 6770 4460 6830 4490
rect 6870 4486 6882 4520
rect 7058 4490 7450 4520
rect 7058 4486 7070 4490
rect 6870 4480 7070 4486
rect 6770 4410 6780 4460
rect 6450 4350 6780 4410
rect 6770 4320 6780 4350
rect 6820 4320 6830 4460
rect 7290 4411 7360 4420
rect 7290 4410 7299 4411
rect 6980 4408 7299 4410
rect 6870 4402 7299 4408
rect 6870 4368 6882 4402
rect 7058 4368 7299 4402
rect 6870 4362 7299 4368
rect 6980 4360 7299 4362
rect 7290 4359 7299 4360
rect 7351 4359 7360 4411
rect 7290 4350 7360 4359
rect 6770 4290 6830 4320
rect 6870 4284 7070 4290
rect 6870 4250 6882 4284
rect 7058 4280 7070 4284
rect 7400 4280 7450 4490
rect 7058 4250 7450 4280
rect 6870 4244 7450 4250
rect 6980 4230 7450 4244
rect 7540 4100 7590 5000
rect 7710 4410 7770 7150
rect 8030 5130 8090 7250
rect 8390 5466 8442 5472
rect 8390 5408 8442 5414
rect 8391 5180 8441 5408
rect 8540 5180 8600 5200
rect 8270 5166 8550 5180
rect 8170 5160 8550 5166
rect 8030 5100 8130 5130
rect 8170 5126 8182 5160
rect 8358 5130 8550 5160
rect 8590 5130 8600 5180
rect 8358 5126 8370 5130
rect 8170 5120 8370 5126
rect 8540 5110 8600 5130
rect 8030 4960 8080 5100
rect 8120 4960 8130 5100
rect 8270 5048 8880 5050
rect 8170 5042 8880 5048
rect 8170 5008 8182 5042
rect 8358 5008 8880 5042
rect 8170 5002 8880 5008
rect 8270 5000 8880 5002
rect 8030 4930 8130 4960
rect 8550 4930 8610 4950
rect 8170 4924 8560 4930
rect 8170 4890 8182 4924
rect 8358 4890 8560 4924
rect 8170 4884 8560 4890
rect 8270 4880 8560 4884
rect 8600 4880 8610 4930
rect 8448 4540 8512 4880
rect 8550 4860 8610 4880
rect 8290 4526 8750 4540
rect 8170 4520 8750 4526
rect 8070 4460 8130 4490
rect 8170 4486 8182 4520
rect 8358 4490 8750 4520
rect 8358 4486 8370 4490
rect 8170 4480 8370 4486
rect 8070 4410 8080 4460
rect 7710 4350 8080 4410
rect 8070 4320 8080 4350
rect 8120 4320 8130 4460
rect 8590 4411 8660 4420
rect 8590 4410 8599 4411
rect 8280 4408 8599 4410
rect 8170 4402 8599 4408
rect 8170 4368 8182 4402
rect 8358 4368 8599 4402
rect 8170 4362 8599 4368
rect 8280 4360 8599 4362
rect 8590 4359 8599 4360
rect 8651 4359 8660 4411
rect 8590 4350 8660 4359
rect 8070 4290 8130 4320
rect 8170 4284 8370 4290
rect 8170 4250 8182 4284
rect 8358 4280 8370 4284
rect 8700 4280 8750 4490
rect 8358 4250 8750 4280
rect 8170 4244 8750 4250
rect 8280 4230 8750 4244
rect 8830 4100 8880 5000
rect 9050 4390 9110 7350
rect 9330 5130 9390 7450
rect 9702 5466 9754 5472
rect 9702 5408 9754 5414
rect 9703 5180 9753 5408
rect 9830 5180 9890 5200
rect 9560 5166 9840 5180
rect 9460 5160 9840 5166
rect 9330 5100 9420 5130
rect 9460 5126 9472 5160
rect 9648 5130 9840 5160
rect 9880 5130 9890 5180
rect 9648 5126 9660 5130
rect 9460 5120 9660 5126
rect 9830 5110 9890 5130
rect 9330 4960 9370 5100
rect 9410 4960 9420 5100
rect 9560 5048 10170 5050
rect 9460 5042 10170 5048
rect 9460 5008 9472 5042
rect 9648 5008 10170 5042
rect 9460 5002 10170 5008
rect 9560 5000 10170 5002
rect 9330 4930 9420 4960
rect 9840 4930 9900 4950
rect 9460 4924 9850 4930
rect 9460 4890 9472 4924
rect 9648 4890 9850 4924
rect 9460 4884 9850 4890
rect 9560 4880 9850 4884
rect 9890 4880 9900 4930
rect 9760 4860 9900 4880
rect 9760 4832 9872 4860
rect 9760 4540 9824 4832
rect 9570 4526 10030 4540
rect 9450 4520 10030 4526
rect 9350 4460 9410 4490
rect 9450 4486 9462 4520
rect 9638 4490 10030 4520
rect 9638 4486 9650 4490
rect 9450 4480 9650 4486
rect 9350 4390 9360 4460
rect 9050 4330 9360 4390
rect 9350 4320 9360 4330
rect 9400 4320 9410 4460
rect 9870 4411 9940 4420
rect 9870 4410 9879 4411
rect 9560 4408 9879 4410
rect 9450 4402 9879 4408
rect 9450 4368 9462 4402
rect 9638 4368 9879 4402
rect 9450 4362 9879 4368
rect 9560 4360 9879 4362
rect 9870 4359 9879 4360
rect 9931 4359 9940 4411
rect 9870 4350 9940 4359
rect 9350 4290 9410 4320
rect 9450 4284 9650 4290
rect 9450 4250 9462 4284
rect 9638 4280 9650 4284
rect 9980 4280 10030 4490
rect 9638 4250 10030 4280
rect 9450 4244 10030 4250
rect 9560 4230 10030 4244
rect 10120 4100 10170 5000
rect -4730 4070 10190 4100
rect -4730 4010 540 4070
rect 600 4010 10190 4070
rect -4730 4000 10190 4010
rect -4730 3906 9960 3930
rect -4730 3896 -3021 3906
rect -5256 3830 -5250 3890
rect -5190 3830 -5184 3890
rect -4730 3844 -4301 3896
rect -4249 3854 -3021 3896
rect -2969 3854 -1721 3906
rect -1669 3854 -441 3906
rect -389 3854 859 3906
rect 911 3854 2139 3906
rect 2191 3854 3439 3906
rect 3491 3854 4719 3906
rect 4771 3854 6019 3906
rect 6071 3854 7299 3906
rect 7351 3854 8599 3906
rect 8651 3854 9879 3906
rect 9931 3854 9960 3906
rect -4249 3844 9960 3854
rect -4730 3830 9960 3844
rect -180 2850 -60 2860
rect -180 2790 -170 2850
rect -70 2790 -60 2850
rect -180 2780 -60 2790
rect -240 2560 -100 2740
rect -20 2700 40 3830
rect 540 3520 600 3526
rect -240 2380 -180 2560
rect 100 2380 160 2760
rect 400 2380 460 2800
rect 540 2700 600 3460
rect 2340 3380 2420 3390
rect 2340 3320 2350 3380
rect 2410 3320 2420 3380
rect 2340 3310 2420 3320
rect 2350 3280 2410 3310
rect 2200 3250 2280 3260
rect 2200 3190 2210 3250
rect 2270 3190 2280 3250
rect 2350 3220 3720 3280
rect 3780 3220 3790 3280
rect 2200 3180 2280 3190
rect 2060 3130 2140 3140
rect 2060 3070 2070 3130
rect 2130 3080 2140 3130
rect 2210 3120 4770 3180
rect 4830 3120 4836 3180
rect 5820 3080 5900 3090
rect 2130 3070 5830 3080
rect 2060 3060 5830 3070
rect 1910 3040 1990 3050
rect 1910 2980 1920 3040
rect 1980 2980 1990 3040
rect 2070 3020 5830 3060
rect 5890 3020 5900 3080
rect 5820 3010 5900 3020
rect 6860 2980 6920 2986
rect 1910 2970 6860 2980
rect 1920 2920 6860 2970
rect 6860 2914 6920 2920
rect 7910 2890 7970 2896
rect 1744 2830 1750 2890
rect 1810 2880 6830 2890
rect 6950 2880 7910 2890
rect 1810 2830 7910 2880
rect 7910 2824 7970 2830
rect 8339 2893 8429 2899
rect 680 2620 820 2800
rect 8339 2790 8429 2803
rect 4160 2720 8430 2790
rect 580 2560 730 2580
rect 580 2480 600 2560
rect 710 2520 730 2560
rect 700 2480 730 2520
rect 580 2470 730 2480
rect 760 2380 820 2620
rect -240 2370 820 2380
rect -240 2320 240 2370
rect 230 2290 240 2320
rect 320 2320 820 2370
rect 320 2290 330 2320
rect 230 2280 330 2290
rect 7904 2196 7976 2202
rect -2540 2140 -2460 2146
rect 3708 2124 3714 2196
rect 3786 2124 3792 2196
rect 4758 2124 4764 2196
rect 4836 2124 4842 2196
rect 5818 2124 5824 2196
rect 5896 2124 5902 2196
rect 6848 2124 6854 2196
rect 6926 2124 6932 2196
rect 7898 2136 7904 2196
rect 7976 2136 7982 2196
rect 7898 2130 7910 2136
rect 7970 2130 7982 2136
rect 7898 2124 7982 2130
rect -3586 1920 -3580 2000
rect -3500 1920 -3494 2000
rect -3580 1820 -3500 1920
rect -2540 1840 -2460 2060
rect -380 2010 -180 2040
rect -470 2000 -350 2010
rect -1500 1920 -350 2000
rect -1500 1840 -1420 1920
rect -470 1870 -350 1920
rect -210 1870 -180 2010
rect -460 1840 -180 1870
rect -10200 1800 -9600 1806
rect -9600 1750 -4100 1800
rect -9600 1500 -4350 1750
rect -4200 1500 -4100 1750
rect 4150 1570 4250 1670
rect -9600 1200 -4100 1500
rect 4154 1446 4245 1570
rect 5210 1450 5290 1590
rect 4148 1355 4154 1446
rect 4245 1355 4251 1446
rect 5190 1430 5310 1450
rect 5190 1350 5210 1430
rect 5290 1350 5310 1430
rect 5190 1330 5310 1350
rect -4020 1300 -3920 1320
rect -4020 1240 -4000 1300
rect -3940 1240 -3920 1300
rect -4020 1220 -3920 1240
rect -3000 1300 -2900 1320
rect -3000 1240 -2980 1300
rect -2920 1240 -2900 1300
rect -3000 1220 -2900 1240
rect -1940 1300 -1840 1320
rect -1940 1240 -1920 1300
rect -1860 1240 -1840 1300
rect -1940 1220 -1840 1240
rect -920 1300 -820 1320
rect -920 1240 -900 1300
rect -840 1240 -820 1300
rect -920 1220 -820 1240
rect -10200 1194 -9600 1200
rect 379 796 501 802
rect -3580 620 -2440 680
rect -4065 549 -3755 561
rect -10225 525 -9575 531
rect -5300 525 -4140 540
rect -9575 400 -4140 525
rect -4065 400 -4059 549
rect -9575 365 -4059 400
rect -9575 55 -5065 365
rect -4755 251 -4059 365
rect -3761 400 -3755 549
rect -3761 251 -3750 400
rect -4755 55 -3750 251
rect -2520 180 -2440 620
rect -1500 380 -1420 680
rect -1320 380 -1240 386
rect -1660 340 -1580 346
rect -1500 300 -1320 380
rect -1320 294 -1240 300
rect -1660 240 -1580 260
rect -460 240 -380 680
rect 379 668 501 674
rect -2890 170 -2790 176
rect -2790 70 -2750 170
rect -2520 80 -2290 180
rect -2190 160 -2184 180
rect -1660 160 -380 240
rect 6265 475 6335 1635
rect 7270 1565 7380 1670
rect 8960 1640 9060 2180
rect 9415 2095 9515 2185
rect 9605 2095 9611 2185
rect 7265 1480 7380 1565
rect 8350 1550 9060 1640
rect 6265 405 7115 475
rect 4409 165 4415 235
rect 4485 165 4491 235
rect -2190 90 -1820 160
rect -2190 80 -2184 90
rect -2890 64 -2760 70
rect -9575 50 -3750 55
rect -9575 -120 -4140 50
rect -2830 10 -2760 64
rect -2830 -60 -2450 10
rect -1890 -20 -1820 90
rect 500 35 2250 50
rect 500 -55 650 35
rect 740 0 2250 35
rect 2509 25 2515 95
rect 2585 25 2880 95
rect 740 -55 750 0
rect 2810 -50 2880 25
rect -9575 -125 -5275 -120
rect -10225 -131 -9575 -125
rect -4000 -1480 -3920 -1160
rect 120 -1460 460 -1400
rect -4000 -2180 -3880 -1480
rect -392 -1580 -234 -1518
rect 120 -1580 180 -1460
rect -392 -1660 -300 -1580
rect -220 -1660 180 -1580
rect -392 -1686 -234 -1660
rect 100 -1760 200 -1750
rect 100 -1800 120 -1760
rect 180 -1800 200 -1760
rect 100 -1810 200 -1800
rect -4000 -2300 -3500 -2180
rect -3620 -4100 -3500 -2300
rect 130 -3560 170 -1810
rect 260 -1820 320 -1620
rect 400 -1660 460 -1460
rect 500 -1820 550 -55
rect 640 -60 750 -55
rect 260 -1850 550 -1820
rect 660 -1780 780 -1140
rect 4415 -1580 4485 165
rect 6265 80 6335 405
rect 6875 235 6945 241
rect 6210 -60 6360 80
rect 6875 -10 6945 165
rect 7045 185 7115 405
rect 7265 365 7355 1480
rect 8780 1050 8880 1550
rect 8780 950 8970 1050
rect 9070 950 9076 1050
rect 8198 760 8402 766
rect 8850 760 9070 780
rect 8198 580 8210 760
rect 8390 580 8870 760
rect 9050 580 9070 760
rect 8198 574 8402 580
rect 8850 560 9070 580
rect 7259 275 7265 365
rect 7355 275 7361 365
rect 7045 115 7275 185
rect 7205 65 7275 115
rect 7205 -5 8775 65
rect 6860 -20 6945 -10
rect 6875 -65 6945 -20
rect 4250 -1650 4485 -1580
rect 4640 -1640 4800 -1160
rect 260 -1880 500 -1850
rect 660 -1900 860 -1780
rect 980 -1900 986 -1780
rect 4634 -1800 4640 -1640
rect 4800 -1800 4806 -1640
rect 8705 -2935 8775 -5
rect 9400 -2534 9560 -2520
rect 9400 -2666 9414 -2534
rect 9546 -2666 9560 -2534
rect 9400 -2680 9560 -2666
rect 8705 -3005 13760 -2935
rect 7030 -3110 7170 -3104
rect 7170 -3114 7330 -3110
rect 7170 -3120 7332 -3114
rect 8890 -3120 9010 -3110
rect 13500 -3120 13560 -3114
rect 7170 -3220 7220 -3120
rect 7320 -3220 8900 -3120
rect 9000 -3220 9010 -3120
rect 7170 -3226 7332 -3220
rect 7170 -3250 7330 -3226
rect 8890 -3230 9010 -3220
rect 11920 -3180 13500 -3120
rect 7030 -3256 7170 -3250
rect 5334 -3554 5386 -3548
rect 130 -3600 5334 -3560
rect 5334 -3612 5386 -3606
rect 4440 -3830 4540 -3824
rect -96 -3930 -90 -3830
rect 10 -3930 4440 -3830
rect 11920 -3840 11980 -3180
rect 13500 -3186 13560 -3180
rect 13690 -3230 13760 -3005
rect 12890 -3290 14020 -3230
rect 12400 -3820 12480 -3800
rect 4440 -3936 4540 -3930
rect 5150 -3900 11990 -3840
rect 12400 -3900 12420 -3820
rect 12460 -3900 12480 -3820
rect 13488 -3876 13494 -3804
rect 13566 -3876 13572 -3804
rect -10850 -4200 -9950 -4194
rect -9950 -5100 -6050 -4200
rect -3620 -4226 -3500 -4220
rect 3960 -4100 4080 -4094
rect 3960 -4400 4080 -4220
rect 5150 -4550 5210 -3900
rect 12400 -3920 12480 -3900
rect 11080 -4090 11300 -4070
rect 8184 -4204 8296 -4198
rect 8184 -4210 8196 -4204
rect 8184 -4310 8190 -4210
rect 8184 -4316 8196 -4310
rect 8296 -4316 8302 -4204
rect 11080 -4270 11100 -4090
rect 11280 -4270 11300 -4090
rect 11080 -4290 11300 -4270
rect 8184 -4322 8296 -4316
rect 11540 -4320 11560 -4200
rect 11674 -4320 11700 -4200
rect 11540 -4340 11700 -4320
rect 5150 -4616 5210 -4610
rect 8100 -4500 12970 -4400
rect 13940 -4450 14020 -4430
rect 13940 -4500 14340 -4450
rect 3694 -4780 3700 -4660
rect 3820 -4780 3826 -4660
rect 8100 -4690 8200 -4500
rect -10850 -5106 -9950 -5100
rect -6950 -5350 -6050 -5100
rect -4000 -5350 -3760 -4840
rect 3700 -4900 3820 -4780
rect 4434 -4790 4440 -4690
rect 4540 -4790 8200 -4690
rect 8290 -4650 10030 -4590
rect 7320 -4824 7420 -4790
rect 7308 -4830 7432 -4824
rect 4040 -5080 4640 -4920
rect 4800 -5080 4806 -4920
rect 7308 -4930 7320 -4830
rect 7420 -4930 7432 -4830
rect 7308 -4936 7432 -4930
rect -6950 -6300 -3760 -5350
rect 5960 -5404 6140 -5400
rect 5960 -5556 5974 -5404
rect 6126 -5556 6140 -5404
rect 5960 -5560 6140 -5556
rect 4100 -5810 4250 -5800
rect 4100 -5890 4110 -5810
rect 4240 -5890 4250 -5810
rect 4100 -5900 4250 -5890
rect 3850 -6110 4000 -6100
rect 3850 -6190 3860 -6110
rect 3990 -6190 4000 -6110
rect 3850 -6200 4000 -6190
rect 4560 -6200 4640 -6120
rect -6950 -6350 -6050 -6300
rect -4000 -6600 -3760 -6300
rect 4320 -6220 4640 -6200
rect 5100 -6220 5160 -6120
rect 5600 -6220 5660 -6120
rect 6120 -6220 6180 -6120
rect 6640 -6220 6700 -6120
rect 7160 -6220 7220 -6120
rect 4320 -6280 7960 -6220
rect 4320 -6340 4400 -6280
rect 4200 -6420 4400 -6340
rect 8020 -6460 8080 -5980
rect 7420 -6520 8080 -6460
rect 4640 -6580 7480 -6520
rect 4840 -6740 4900 -6580
rect 5340 -6740 5400 -6580
rect 5860 -6740 5920 -6580
rect 6380 -6740 6440 -6580
rect 6900 -6740 6960 -6580
rect 7420 -6740 7480 -6580
rect 7800 -6780 7860 -6520
rect 7800 -6820 7880 -6780
rect 8290 -6900 8350 -4650
rect 9970 -4750 10030 -4650
rect 10584 -4690 10590 -4590
rect 10690 -4690 10696 -4590
rect 14280 -4650 14340 -4500
rect 14564 -4560 14570 -4480
rect 14650 -4560 14656 -4480
rect 14269 -4655 14275 -4650
rect 10590 -4750 10690 -4690
rect 13950 -4695 14020 -4690
rect 14105 -4695 14275 -4655
rect 13950 -4700 14275 -4695
rect 13940 -4720 14275 -4700
rect 14345 -4720 14370 -4650
rect 13940 -4725 14345 -4720
rect 13940 -4765 14175 -4725
rect 14570 -4740 14650 -4560
rect 13940 -4770 14020 -4765
rect 12050 -6390 12130 -5850
rect 12020 -6440 12160 -6390
rect 12014 -6580 12020 -6440
rect 12160 -6580 12166 -6440
rect 16025 -6515 16135 -5965
rect 16025 -6631 16135 -6625
rect 8020 -6960 8350 -6900
rect 8020 -7000 8240 -6960
rect 8160 -7200 8240 -7000
rect 8160 -7280 9080 -7200
rect 8160 -7340 8240 -7280
rect 7840 -7360 8240 -7340
rect 5150 -7430 5210 -7424
rect 5328 -7486 5334 -7434
rect 5386 -7486 5392 -7434
rect 5150 -13410 5210 -7490
rect 5340 -13180 5380 -7486
rect 7840 -7500 7860 -7360
rect 8220 -7500 8240 -7360
rect 8780 -7380 8840 -7280
rect 9020 -7380 9080 -7280
rect 9320 -7280 9660 -7220
rect 9320 -7330 9390 -7280
rect 7840 -7520 8240 -7500
rect 8900 -7620 8960 -7480
rect 9270 -7540 9390 -7330
rect 9590 -7360 9660 -7280
rect 11580 -7375 11770 -7360
rect 8754 -7680 8760 -7620
rect 8820 -7680 8960 -7620
rect 9000 -7580 9100 -7570
rect 9270 -7580 9350 -7540
rect 9000 -7620 9020 -7580
rect 9080 -7620 9100 -7580
rect 9000 -7630 9100 -7620
rect 9250 -7600 9350 -7580
rect 9020 -10710 9080 -7630
rect 9250 -7670 9260 -7600
rect 9340 -7670 9350 -7600
rect 9470 -7660 9520 -7500
rect 11580 -7525 11600 -7375
rect 11750 -7525 11770 -7375
rect 11580 -7540 11770 -7525
rect 9590 -7580 9670 -7570
rect 9590 -7620 9610 -7580
rect 9650 -7620 9670 -7580
rect 9590 -7630 9670 -7620
rect 9250 -7680 9350 -7670
rect 9450 -7670 9540 -7660
rect 9450 -7730 9460 -7670
rect 9530 -7730 9540 -7670
rect 9450 -7740 9540 -7730
rect 9600 -10550 9660 -7630
rect 11695 -7775 11805 -7769
rect 11805 -7885 12275 -7775
rect 12385 -7885 12391 -7775
rect 11695 -7891 11805 -7885
rect 9600 -10610 16090 -10550
rect 9020 -10770 15090 -10710
rect 14448 -13180 14454 -13174
rect 5340 -13220 14454 -13180
rect 14448 -13226 14454 -13220
rect 14506 -13226 14512 -13174
rect 5150 -13476 5210 -13470
rect 15030 -13820 15090 -10770
rect 15030 -13886 15090 -13880
rect 16030 -13820 16090 -10610
rect 16030 -13886 16090 -13880
<< via1 >>
rect -7810 6830 -7750 6890
rect -7690 6710 -7630 6770
rect -7570 6590 -7510 6650
rect -7470 6490 -7410 6550
rect -7350 6390 -7290 6450
rect -7230 6290 -7170 6350
rect -7090 6190 -7030 6250
rect -6970 6090 -6910 6150
rect -6850 5990 -6790 6050
rect -6730 5890 -6670 5950
rect -6590 5790 -6530 5850
rect -6470 5690 -6410 5750
rect -6350 5590 -6290 5650
rect -6250 5450 -6190 5510
rect -6130 5330 -6070 5390
rect -6010 5230 -5950 5290
rect -5910 5130 -5850 5190
rect -5790 5030 -5730 5090
rect -5690 4910 -5630 4970
rect -5590 4810 -5530 4870
rect -4486 5129 -4434 5181
rect -5250 4990 -5190 5050
rect -5470 4710 -5410 4770
rect -4301 4359 -4249 4411
rect -3210 5254 -3158 5306
rect -3021 4359 -2969 4411
rect -1930 5430 -1878 5482
rect -1721 4359 -1669 4411
rect -650 5542 -598 5594
rect -441 4359 -389 4411
rect 646 5350 698 5402
rect 859 4359 911 4411
rect 1926 5510 1978 5562
rect 2139 4359 2191 4411
rect 3238 5686 3290 5738
rect 3439 4359 3491 4411
rect 4534 5926 4586 5978
rect 4176 5376 4240 5440
rect 4719 4359 4771 4411
rect 5814 6134 5866 6186
rect 6019 4359 6071 4411
rect 7110 5414 7162 5466
rect 7299 4359 7351 4411
rect 8390 5414 8442 5466
rect 8599 4359 8651 4411
rect 9702 5414 9754 5466
rect 9879 4359 9931 4411
rect 540 4010 600 4070
rect -5250 3830 -5190 3890
rect -4301 3844 -4249 3896
rect -3021 3854 -2969 3906
rect -1721 3854 -1669 3906
rect -441 3854 -389 3906
rect 859 3854 911 3906
rect 2139 3854 2191 3906
rect 3439 3854 3491 3906
rect 4719 3854 4771 3906
rect 6019 3854 6071 3906
rect 7299 3854 7351 3906
rect 8599 3854 8651 3906
rect 9879 3854 9931 3906
rect -170 2840 -70 2850
rect -170 2800 -160 2840
rect -160 2800 -80 2840
rect -80 2800 -70 2840
rect -170 2790 -70 2800
rect 540 3460 600 3520
rect 2350 3320 2410 3380
rect 2210 3190 2270 3250
rect 3720 3220 3780 3280
rect 2070 3070 2130 3130
rect 4770 3120 4830 3180
rect 1920 2980 1980 3040
rect 5830 3020 5890 3080
rect 6860 2920 6920 2980
rect 1750 2830 1810 2890
rect 7910 2830 7970 2890
rect 8339 2803 8429 2893
rect 600 2520 700 2560
rect 600 2480 700 2520
rect 240 2290 320 2370
rect -2540 2060 -2460 2140
rect 3714 2190 3786 2196
rect 3714 2130 3720 2190
rect 3720 2130 3780 2190
rect 3780 2130 3786 2190
rect 3714 2124 3786 2130
rect 4764 2190 4836 2196
rect 4764 2130 4770 2190
rect 4770 2130 4830 2190
rect 4830 2130 4836 2190
rect 4764 2124 4836 2130
rect 5824 2190 5896 2196
rect 5824 2130 5830 2190
rect 5830 2130 5890 2190
rect 5890 2130 5896 2190
rect 5824 2124 5896 2130
rect 6854 2190 6926 2196
rect 6854 2130 6860 2190
rect 6860 2130 6920 2190
rect 6920 2130 6926 2190
rect 6854 2124 6926 2130
rect 7904 2190 7976 2196
rect 7904 2136 7910 2190
rect 7910 2136 7970 2190
rect 7970 2136 7976 2190
rect -3580 1920 -3500 2000
rect -350 1870 -210 2010
rect -10200 1200 -9600 1800
rect 4154 1355 4245 1446
rect 5210 1350 5290 1430
rect -4000 1240 -3960 1300
rect -3960 1240 -3940 1300
rect -2980 1240 -2920 1300
rect -1920 1240 -1860 1300
rect -900 1240 -840 1300
rect 379 790 501 796
rect 379 680 385 790
rect 385 680 495 790
rect 495 680 501 790
rect -10225 -125 -9575 525
rect -1660 260 -1580 340
rect -1320 300 -1240 380
rect 379 674 501 680
rect -2890 70 -2790 170
rect -2290 80 -2190 180
rect 9515 2095 9605 2185
rect 4415 165 4485 235
rect 650 -55 740 35
rect 2515 25 2585 95
rect -300 -1660 -220 -1580
rect 6875 165 6945 235
rect 8970 950 9070 1050
rect 8870 580 9050 760
rect 7265 275 7355 365
rect 860 -1900 980 -1780
rect 4640 -1800 4800 -1640
rect 9414 -2540 9546 -2534
rect 9414 -2660 9420 -2540
rect 9420 -2660 9540 -2540
rect 9540 -2660 9546 -2540
rect 9414 -2666 9546 -2660
rect 7030 -3250 7170 -3110
rect 8900 -3220 9000 -3120
rect 13500 -3180 13560 -3120
rect 5334 -3606 5386 -3554
rect -90 -3930 10 -3830
rect 4440 -3930 4540 -3830
rect 13494 -3810 13566 -3804
rect 13494 -3870 13500 -3810
rect 13500 -3870 13560 -3810
rect 13560 -3870 13566 -3810
rect 13494 -3876 13566 -3870
rect -10850 -5100 -9950 -4200
rect -3620 -4220 -3500 -4100
rect 3960 -4220 4080 -4100
rect 8196 -4210 8296 -4204
rect 8196 -4310 8290 -4210
rect 8290 -4310 8296 -4210
rect 8196 -4316 8296 -4310
rect 11100 -4096 11280 -4090
rect 11100 -4264 11106 -4096
rect 11106 -4264 11274 -4096
rect 11274 -4264 11280 -4096
rect 11100 -4270 11280 -4264
rect 11560 -4206 11674 -4200
rect 11560 -4314 11566 -4206
rect 11566 -4314 11674 -4206
rect 11560 -4320 11674 -4314
rect 5150 -4610 5210 -4550
rect 3700 -4780 3820 -4660
rect 4440 -4790 4540 -4690
rect 4640 -5080 4800 -4920
rect 5974 -5410 6126 -5404
rect 5974 -5550 5980 -5410
rect 5980 -5550 6120 -5410
rect 6120 -5550 6126 -5410
rect 5974 -5556 6126 -5550
rect 4110 -5890 4240 -5810
rect 3860 -6190 3990 -6110
rect 10590 -4690 10690 -4590
rect 14570 -4560 14650 -4480
rect 14275 -4720 14345 -4650
rect 12020 -6580 12160 -6440
rect 16025 -6625 16135 -6515
rect 5150 -7490 5210 -7430
rect 5334 -7486 5386 -7434
rect 7860 -7500 8220 -7360
rect 8760 -7680 8820 -7620
rect 9260 -7670 9340 -7600
rect 11600 -7381 11750 -7375
rect 11600 -7519 11606 -7381
rect 11606 -7519 11744 -7381
rect 11744 -7519 11750 -7381
rect 11600 -7525 11750 -7519
rect 9460 -7730 9530 -7670
rect 11695 -7885 11805 -7775
rect 12275 -7885 12385 -7775
rect 14454 -13226 14506 -13174
rect 5150 -13470 5210 -13410
rect 15030 -13880 15090 -13820
rect 16030 -13880 16090 -13820
<< metal2 >>
rect -8400 7700 -7600 9200
rect -6700 7700 -5900 9200
rect -5100 7700 -4300 9200
rect -3500 7700 -2700 9200
rect -1900 7700 -1100 9200
rect -300 7700 500 9200
rect 1300 7700 2100 9200
rect 2900 7700 3700 9200
rect 4500 7700 5300 9200
rect 6100 7700 6900 9200
rect 7700 7700 8500 9200
rect 9300 7700 10100 9200
rect -8000 7680 -7880 7700
rect -6400 7680 -6280 7700
rect -4800 7680 -4680 7700
rect -3200 7680 -3080 7700
rect -1600 7680 -1480 7700
rect 0 7680 120 7700
rect 1600 7680 1720 7700
rect 3200 7680 3320 7700
rect 4800 7680 4920 7700
rect 6400 7680 6520 7700
rect 8000 7680 8120 7700
rect -7966 7004 -7906 7680
rect -6366 7196 -6306 7680
rect -4782 7372 -4722 7680
rect -3182 7374 -3122 7680
rect -1566 7580 -1506 7680
rect 34 7644 94 7680
rect 27 7588 36 7644
rect 92 7588 101 7644
rect 1634 7628 1694 7680
rect 3234 7628 3294 7680
rect 34 7586 94 7588
rect -1573 7524 -1564 7580
rect -1508 7524 -1499 7580
rect 1627 7572 1636 7628
rect 1692 7572 1701 7628
rect 3227 7572 3236 7628
rect 3292 7572 3301 7628
rect 4818 7612 4878 7680
rect 6434 7628 6494 7680
rect 8018 7628 8078 7680
rect 1634 7570 1694 7572
rect 3234 7570 3294 7572
rect 4811 7556 4820 7612
rect 4876 7556 4885 7612
rect 6427 7572 6436 7628
rect 6492 7572 6501 7628
rect 8018 7572 8020 7628
rect 8076 7572 8078 7628
rect 9600 7600 9800 7700
rect 9634 7586 9758 7600
rect 6434 7570 6494 7572
rect 8018 7570 8078 7572
rect 8020 7563 8076 7570
rect 4818 7554 4878 7556
rect -1566 7522 -1506 7524
rect 9698 7516 9758 7586
rect 9691 7460 9700 7516
rect 9756 7460 9765 7516
rect 9698 7458 9758 7460
rect -652 7374 -596 7381
rect -3182 7372 -594 7374
rect -4789 7316 -4780 7372
rect -4724 7316 -4715 7372
rect -3182 7316 -652 7372
rect -596 7316 -594 7372
rect -4782 7314 -4722 7316
rect -3182 7314 -594 7316
rect -652 7307 -596 7314
rect -6373 7140 -6364 7196
rect -6308 7140 -6299 7196
rect -6366 7138 -6306 7140
rect -7973 6948 -7964 7004
rect -7908 6948 -7899 7004
rect -7966 6946 -7906 6948
rect -7816 6830 -7810 6890
rect -7750 6830 -7744 6890
rect -11500 1900 -10900 1909
rect -10900 1300 -10200 1800
rect -11500 1200 -10200 1300
rect -9600 1200 -9594 1800
rect -11500 1100 -10900 1200
rect -12500 500 -11900 509
rect -11500 500 -10900 600
rect -10300 500 -10225 525
rect -12600 -100 -12500 500
rect -11900 -100 -10225 500
rect -12500 -109 -11900 -100
rect -11500 -200 -10900 -100
rect -10300 -125 -10225 -100
rect -9575 -125 -9569 525
rect -11500 -4450 -10850 -4200
rect -9950 -5100 -9944 -4200
rect -11500 -5109 -10850 -5100
rect -12200 -6000 -10700 -5600
rect -12200 -6030 -10660 -6000
rect -7810 -6030 -7750 6830
rect -7696 6710 -7690 6770
rect -7630 6710 -7624 6770
rect -12200 -6090 -7750 -6030
rect -12200 -6120 -10660 -6090
rect -12200 -6400 -10700 -6120
rect -12200 -7000 -10700 -6600
rect -12200 -7030 -10660 -7000
rect -7690 -7030 -7630 6710
rect -12200 -7090 -7630 -7030
rect -7570 6650 -7510 6656
rect -12200 -7120 -10660 -7090
rect -12200 -7400 -10700 -7120
rect -12200 -8000 -10700 -7600
rect -12200 -8030 -10660 -8000
rect -7570 -8030 -7510 6590
rect -12200 -8090 -7510 -8030
rect -7470 6550 -7410 6556
rect -12200 -8120 -10670 -8090
rect -12200 -8400 -10700 -8120
rect -7470 -8490 -7410 6490
rect -8270 -8550 -7410 -8490
rect -7350 6450 -7290 6456
rect -12200 -9000 -10700 -8600
rect -12200 -9030 -10660 -9000
rect -8270 -9030 -8210 -8550
rect -7350 -8590 -7290 6390
rect -12200 -9090 -8210 -9030
rect -8170 -8650 -7290 -8590
rect -7230 6350 -7170 6356
rect -12200 -9120 -10660 -9090
rect -12200 -9400 -10700 -9120
rect -12200 -10000 -10700 -9600
rect -12200 -10030 -10660 -10000
rect -8170 -10030 -8110 -8650
rect -7230 -8710 -7170 6290
rect -12200 -10090 -8110 -10030
rect -8050 -8770 -7170 -8710
rect -7090 6250 -7030 6256
rect -12200 -10120 -10660 -10090
rect -12200 -10400 -10700 -10120
rect -12200 -11000 -10700 -10600
rect -12200 -11030 -10660 -11000
rect -8050 -11030 -7990 -8770
rect -7090 -8830 -7030 6190
rect 5792 6190 5888 6208
rect -12200 -11090 -7990 -11030
rect -7910 -8890 -7030 -8830
rect -6970 6150 -6910 6156
rect 5792 6130 5810 6190
rect 5870 6130 5888 6190
rect 5792 6112 5888 6130
rect -12200 -11120 -10660 -11090
rect -12200 -11400 -10700 -11120
rect -12200 -12000 -10700 -11600
rect -12200 -12030 -10660 -12000
rect -7910 -12030 -7850 -8890
rect -6970 -8990 -6910 6090
rect -12200 -12090 -7850 -12030
rect -7790 -9050 -6910 -8990
rect -6850 6050 -6790 6056
rect -12200 -12120 -10660 -12090
rect -12200 -12400 -10700 -12120
rect -7790 -12330 -7730 -9050
rect -6850 -9130 -6790 5990
rect 4512 5982 4608 6000
rect -10150 -12390 -7730 -12330
rect -7650 -9190 -6790 -9130
rect -6730 5950 -6670 5956
rect -5036 5920 -4980 5925
rect 4512 5922 4530 5982
rect 4590 5922 4608 5982
rect -12200 -13000 -10700 -12600
rect -12200 -13030 -10660 -13000
rect -10150 -13030 -10090 -12390
rect -7650 -12430 -7590 -9190
rect -6730 -9250 -6670 5890
rect -5040 5916 4240 5920
rect -5040 5860 -5036 5916
rect -4980 5860 4240 5916
rect 4512 5904 4608 5922
rect -5040 5856 4240 5860
rect -12200 -13090 -10090 -13030
rect -9970 -12490 -7590 -12430
rect -7550 -9310 -6670 -9250
rect -6590 5850 -6530 5856
rect -5036 5851 -4980 5856
rect -12200 -13120 -10660 -13090
rect -12200 -13400 -10700 -13120
rect -10960 -13520 -10400 -13456
rect -10336 -13520 -10327 -13456
rect -10960 -13680 -10896 -13520
rect -9970 -13660 -9910 -12490
rect -7550 -12530 -7490 -9310
rect -6590 -9350 -6530 5790
rect -8970 -12590 -7490 -12530
rect -7430 -9410 -6530 -9350
rect -6470 5750 -6410 5756
rect -8970 -13660 -8910 -12590
rect -7430 -12650 -7370 -9410
rect -6470 -9450 -6410 5690
rect 3216 5742 3312 5760
rect 3216 5682 3234 5742
rect 3294 5682 3312 5742
rect 3216 5664 3312 5682
rect -7970 -12710 -7370 -12650
rect -6970 -9510 -6410 -9450
rect -6350 5650 -6290 5656
rect -6350 -9450 -6290 5590
rect -672 5600 -576 5616
rect -672 5538 -654 5600
rect -594 5538 -576 5600
rect -672 5520 -576 5538
rect 1904 5566 2000 5584
rect -6256 5450 -6250 5510
rect -6190 5450 -6184 5510
rect 1904 5506 1922 5566
rect 1982 5506 2000 5566
rect -1952 5486 -1856 5504
rect 1904 5488 2000 5506
rect -6250 -9330 -6190 5450
rect -1952 5426 -1934 5486
rect -1874 5426 -1856 5486
rect -1952 5424 -1856 5426
rect 4176 5440 4240 5856
rect 646 5406 698 5408
rect -6130 5390 -6070 5396
rect 633 5346 642 5406
rect 702 5346 711 5406
rect 7088 5470 7184 5488
rect 7088 5410 7106 5470
rect 7166 5410 7184 5470
rect 7088 5392 7184 5410
rect 8368 5470 8464 5488
rect 8368 5410 8386 5470
rect 8446 5410 8464 5470
rect 9689 5410 9698 5470
rect 9758 5410 9767 5470
rect 8368 5392 8464 5410
rect 4176 5370 4240 5376
rect 646 5344 698 5346
rect -6130 -9230 -6070 5330
rect -3232 5310 -3136 5328
rect -6010 5290 -5950 5296
rect -6010 -9130 -5950 5230
rect -4490 5250 -4430 5259
rect -5910 5190 -5850 5196
rect -3232 5250 -3214 5310
rect -3154 5250 -3136 5310
rect -3232 5216 -3136 5250
rect -4490 5181 -4430 5190
rect -5910 -9030 -5850 5130
rect -4492 5129 -4486 5181
rect -4434 5129 -4428 5181
rect -5790 5090 -5730 5096
rect -5790 -8930 -5730 5030
rect -5256 4990 -5250 5050
rect -5190 4990 -5184 5050
rect -5690 4970 -5630 4976
rect -5690 -8810 -5630 4910
rect -5590 4870 -5530 4876
rect -5590 -8710 -5530 4810
rect -5470 4770 -5410 4776
rect -5470 -8590 -5410 4710
rect -5250 4610 -5190 4990
rect -5370 4550 -5190 4610
rect -5370 -8490 -5310 4550
rect -4310 4411 -4240 4420
rect -4310 4359 -4301 4411
rect -4249 4359 -4240 4411
rect -4310 4350 -4240 4359
rect -3030 4411 -2960 4420
rect -3030 4359 -3021 4411
rect -2969 4359 -2960 4411
rect -3030 4350 -2960 4359
rect -1730 4411 -1660 4420
rect -1730 4359 -1721 4411
rect -1669 4359 -1660 4411
rect -1730 4350 -1660 4359
rect -450 4411 -380 4420
rect -450 4359 -441 4411
rect -389 4359 -380 4411
rect -450 4350 -380 4359
rect 850 4411 920 4420
rect 850 4359 859 4411
rect 911 4359 920 4411
rect 850 4350 920 4359
rect 2130 4411 2200 4420
rect 2130 4359 2139 4411
rect 2191 4359 2200 4411
rect 2130 4350 2200 4359
rect 3430 4411 3500 4420
rect 3430 4359 3439 4411
rect 3491 4359 3500 4411
rect 3430 4350 3500 4359
rect 4710 4411 4780 4420
rect 4710 4359 4719 4411
rect 4771 4359 4780 4411
rect 4710 4350 4780 4359
rect 6010 4411 6080 4420
rect 6010 4359 6019 4411
rect 6071 4359 6080 4411
rect 6010 4350 6080 4359
rect 7290 4411 7360 4420
rect 7290 4359 7299 4411
rect 7351 4359 7360 4411
rect 7290 4350 7360 4359
rect 8590 4411 8660 4420
rect 8590 4359 8599 4411
rect 8651 4359 8660 4411
rect 8590 4350 8660 4359
rect 9870 4411 9940 4420
rect 9870 4359 9879 4411
rect 9931 4359 9940 4411
rect 9870 4350 9940 4359
rect -4300 3902 -4250 4350
rect -3020 3912 -2970 4350
rect -1720 3912 -1670 4350
rect -440 3912 -390 4350
rect 540 4070 600 4076
rect -3021 3906 -2969 3912
rect -4301 3896 -4249 3902
rect -5250 3890 -5190 3896
rect -3021 3848 -2969 3854
rect -1721 3906 -1669 3912
rect -1721 3848 -1669 3854
rect -441 3906 -389 3912
rect -441 3848 -389 3854
rect -4301 3838 -4249 3844
rect -5250 -8370 -5190 3830
rect -5160 3740 -5100 3749
rect -5160 -8260 -5100 3680
rect -5060 3600 -5000 3609
rect -5060 -8160 -5000 3540
rect 540 3520 600 4010
rect 860 3912 910 4350
rect 859 3906 911 3912
rect 2140 3906 2190 4350
rect 3440 3912 3490 4350
rect 4720 3912 4770 4350
rect 6020 3912 6070 4350
rect 3439 3906 3491 3912
rect 2133 3854 2139 3906
rect 2191 3854 2197 3906
rect 859 3848 911 3854
rect 3439 3848 3491 3854
rect 4719 3906 4771 3912
rect 4719 3848 4771 3854
rect 6019 3906 6071 3912
rect 7300 3906 7350 4350
rect 8600 3912 8650 4350
rect 9880 3912 9930 4350
rect 8599 3906 8651 3912
rect 7293 3854 7299 3906
rect 7351 3854 7357 3906
rect 6019 3848 6071 3854
rect 8599 3848 8651 3854
rect 9879 3906 9931 3912
rect 9879 3848 9931 3854
rect -4960 3460 -4900 3469
rect 534 3460 540 3520
rect 600 3460 606 3520
rect -4960 -8060 -4900 3400
rect 2340 3380 2420 3390
rect -4860 3330 -4800 3339
rect 2340 3320 2350 3380
rect 2410 3320 2420 3380
rect 2340 3310 2420 3320
rect -4860 -7960 -4800 3270
rect 3720 3280 3780 3286
rect 2200 3250 2280 3260
rect -4760 3190 -4700 3199
rect 2200 3190 2210 3250
rect 2270 3190 2280 3250
rect 2200 3180 2280 3190
rect -4760 -7860 -4700 3130
rect 2060 3130 2140 3140
rect 2060 3070 2070 3130
rect 2130 3070 2140 3130
rect 2060 3060 2140 3070
rect 1910 3040 1990 3050
rect 1910 2980 1920 3040
rect 1980 2980 1990 3040
rect 1910 2970 1990 2980
rect 1750 2890 1810 2899
rect -180 2850 -60 2860
rect -430 2840 -170 2850
rect -4660 2790 -170 2840
rect -70 2790 -60 2850
rect 1750 2821 1810 2830
rect -4660 2780 -370 2790
rect -180 2780 -60 2790
rect -4660 -7760 -4600 2780
rect 580 2560 730 2580
rect -4560 2550 -350 2560
rect 580 2550 600 2560
rect -4560 2500 600 2550
rect -4560 -7660 -4500 2500
rect -430 2490 600 2500
rect 580 2480 600 2490
rect 700 2480 730 2560
rect 580 2470 730 2480
rect 230 2370 330 2380
rect 230 2290 240 2370
rect 320 2290 330 2370
rect -2560 2140 -2440 2160
rect -4460 2060 -2920 2120
rect -4460 -7560 -4400 2060
rect -3600 2000 -3480 2020
rect -3600 1920 -3580 2000
rect -3500 1920 -3480 2000
rect -3600 1900 -3480 1920
rect -2980 1980 -2920 2060
rect -2560 2060 -2540 2140
rect -2460 2060 -2440 2140
rect -2560 2040 -2440 2060
rect -380 2010 -180 2040
rect -2980 1920 -840 1980
rect -2980 1320 -2920 1920
rect -900 1320 -840 1920
rect -380 1870 -350 2010
rect -210 1870 -180 2010
rect -380 1840 -180 1870
rect -4020 1300 -3920 1320
rect -4360 1240 -4000 1300
rect -3940 1240 -3920 1300
rect -4360 -7460 -4300 1240
rect -4020 1220 -3920 1240
rect -3000 1300 -2900 1320
rect -3000 1240 -2980 1300
rect -2920 1240 -2900 1300
rect -3000 1220 -2900 1240
rect -1940 1300 -1840 1320
rect -1940 1240 -1920 1300
rect -1860 1240 -1840 1300
rect -1940 1220 -1840 1240
rect -920 1300 -820 1320
rect -920 1240 -900 1300
rect -840 1240 -820 1300
rect -920 1220 -820 1240
rect -4000 540 -3940 1220
rect -1920 540 -1860 1220
rect -4000 480 -1860 540
rect -1340 380 -1220 400
rect -1680 340 -1560 360
rect -1680 260 -1660 340
rect -1580 260 -1560 340
rect -1340 300 -1320 380
rect -1240 300 -1220 380
rect -1340 280 -1220 300
rect -1680 240 -1560 260
rect -2290 180 -2190 186
rect 230 180 330 2290
rect 3720 2210 3780 3220
rect 4770 3180 4830 3186
rect 4770 2210 4830 3120
rect 5820 3080 5900 3090
rect 5820 3020 5830 3080
rect 5890 3020 5900 3080
rect 5820 3010 5900 3020
rect 5830 2210 5890 3010
rect 6854 2920 6860 2980
rect 6920 2920 6926 2980
rect 6860 2210 6920 2920
rect 7904 2830 7910 2890
rect 7970 2830 7976 2890
rect 3700 2196 3800 2210
rect 3700 2124 3714 2196
rect 3786 2124 3800 2196
rect 3700 2110 3800 2124
rect 4750 2196 4850 2210
rect 4750 2124 4764 2196
rect 4836 2124 4850 2196
rect 4750 2110 4850 2124
rect 5810 2196 5910 2210
rect 5810 2124 5824 2196
rect 5896 2124 5910 2196
rect 5810 2110 5910 2124
rect 6840 2196 6940 2210
rect 7910 2196 7970 2830
rect 8333 2803 8339 2893
rect 8429 2803 10493 2893
rect 6840 2124 6854 2196
rect 6926 2124 6940 2196
rect 7898 2136 7904 2196
rect 7976 2136 7982 2196
rect 9515 2185 9605 2191
rect 6840 2110 6940 2124
rect 9515 1520 9605 2095
rect 4140 1446 4260 1460
rect 4140 1355 4154 1446
rect 4245 1355 4260 1446
rect 4140 1340 4260 1355
rect 5190 1430 5310 1450
rect 5190 1350 5210 1430
rect 5290 1350 5310 1430
rect 9515 1405 9600 1520
rect 5190 1330 5310 1350
rect 8665 1315 9600 1405
rect 10403 1405 10493 2803
rect 15700 1405 17200 1800
rect 10403 1315 17200 1405
rect 360 796 520 810
rect 360 674 379 796
rect 501 674 520 796
rect 360 660 520 674
rect 7240 365 7370 380
rect 7240 275 7265 365
rect 7355 275 7370 365
rect 7240 260 7370 275
rect -2896 70 -2890 170
rect -2790 70 -2784 170
rect -2190 80 330 180
rect 4415 235 4485 241
rect 4485 165 6875 235
rect 6945 165 6951 235
rect 4415 159 4485 165
rect 2500 95 2600 110
rect -2290 74 -2190 80
rect 640 35 750 50
rect 640 -55 650 35
rect 740 -55 750 35
rect 2500 25 2515 95
rect 2585 25 2600 95
rect 2500 10 2600 25
rect 640 -60 750 -55
rect -90 -80 10 -71
rect -392 -1550 -234 -1518
rect -392 -1580 -200 -1550
rect -392 -1660 -300 -1580
rect -220 -1660 -200 -1580
rect -392 -1680 -200 -1660
rect -392 -1686 -234 -1680
rect -90 -3830 10 -180
rect 8665 -1570 8755 1315
rect 8970 1050 9070 1056
rect 9070 950 10670 1050
rect 15700 1000 17200 1315
rect 8970 944 9070 950
rect 8850 760 9070 780
rect 8850 580 8870 760
rect 9050 580 9070 760
rect 8850 560 9070 580
rect 10570 130 10670 950
rect 15600 130 17200 400
rect 10570 30 17200 130
rect 15600 -400 17200 30
rect 4640 -1640 4800 -1634
rect 860 -1780 980 -1774
rect 860 -2780 980 -1900
rect 8330 -1660 8755 -1570
rect 860 -2900 4080 -2780
rect -90 -3936 10 -3930
rect 3960 -4100 4080 -2900
rect 4434 -3930 4440 -3830
rect 4540 -3930 4546 -3830
rect -3626 -4220 -3620 -4100
rect -3500 -4220 3820 -4100
rect 3954 -4220 3960 -4100
rect 4080 -4220 4086 -4100
rect 3700 -4660 3820 -4220
rect 3700 -4786 3820 -4780
rect 4440 -4690 4540 -3930
rect 4440 -4796 4540 -4790
rect 4640 -4920 4800 -1800
rect 9400 -2534 9560 -2520
rect 9400 -2666 9414 -2534
rect 9546 -2540 9560 -2534
rect 9546 -2660 11680 -2540
rect 9546 -2666 9560 -2660
rect 9400 -2680 9560 -2666
rect 5980 -3250 7030 -3110
rect 7170 -3250 7176 -3110
rect 8890 -3120 9010 -3110
rect 8890 -3220 8900 -3120
rect 9000 -3220 9010 -3120
rect 8890 -3230 9010 -3220
rect 5328 -3606 5334 -3554
rect 5386 -3606 5392 -3554
rect 5144 -4610 5150 -4550
rect 5210 -4610 5216 -4550
rect 4640 -5086 4800 -5080
rect 4100 -5810 4250 -5800
rect 4100 -5890 4110 -5810
rect 4240 -5890 4250 -5810
rect 4100 -6000 4250 -5890
rect 3850 -6110 4000 -6100
rect 3850 -6190 3860 -6110
rect 3990 -6190 4000 -6110
rect 3850 -6330 4000 -6190
rect -4360 -7520 1940 -7460
rect -4460 -7620 1840 -7560
rect -4560 -7720 1740 -7660
rect -4660 -7820 1640 -7760
rect -4760 -7920 1540 -7860
rect -4860 -8020 1430 -7960
rect -4960 -8120 1330 -8060
rect -5060 -8220 1210 -8160
rect -5160 -8320 1090 -8260
rect -5250 -8430 990 -8370
rect -5370 -8550 870 -8490
rect -5470 -8650 750 -8590
rect -5590 -8770 650 -8710
rect -5690 -8870 90 -8810
rect -5790 -8990 -910 -8930
rect -5910 -9090 -1910 -9030
rect -6010 -9190 -2910 -9130
rect -6130 -9290 -3910 -9230
rect -6250 -9390 -4910 -9330
rect -6350 -9510 -5910 -9450
rect -7970 -13660 -7910 -12710
rect -6970 -13660 -6910 -9510
rect -5970 -13660 -5910 -9510
rect -4970 -13660 -4910 -9390
rect -3970 -13660 -3910 -9290
rect -2970 -13660 -2910 -9190
rect -1970 -13660 -1910 -9090
rect -970 -13660 -910 -8990
rect 30 -13660 90 -8870
rect 590 -13170 650 -8770
rect 690 -13070 750 -8650
rect 810 -12970 870 -8550
rect 930 -12870 990 -8430
rect 1030 -12770 1090 -8320
rect 1150 -12670 1210 -8220
rect 1270 -12570 1330 -8120
rect 1370 -12470 1430 -8020
rect 1480 -12370 1540 -7920
rect 1580 -12270 1640 -7820
rect 1680 -12170 1740 -7720
rect 1780 -12070 1840 -7620
rect 1880 -11970 1940 -7520
rect 3850 -7970 3990 -6330
rect 4135 -7775 4245 -6000
rect 5150 -7430 5210 -4610
rect 5340 -7428 5380 -3606
rect 5980 -5400 6120 -3250
rect 11080 -4090 11300 -4070
rect 8196 -4204 8296 -4198
rect 8296 -4310 10690 -4210
rect 11080 -4270 11100 -4090
rect 11280 -4270 11300 -4090
rect 11560 -4200 11680 -2660
rect 13494 -3180 13500 -3120
rect 13560 -3180 13566 -3120
rect 13500 -3790 13560 -3180
rect 13480 -3804 13580 -3790
rect 13480 -3876 13494 -3804
rect 13566 -3876 13580 -3804
rect 13480 -3890 13580 -3876
rect 11080 -4290 11300 -4270
rect 8196 -4322 8296 -4316
rect 10590 -4590 10690 -4310
rect 11540 -4320 11560 -4200
rect 11674 -4320 11700 -4200
rect 11540 -4340 11700 -4320
rect 14570 -4480 14650 -4474
rect 14570 -4566 14650 -4560
rect 10590 -4696 10690 -4690
rect 14250 -4650 14370 -4630
rect 14250 -4720 14275 -4650
rect 14345 -4720 14370 -4650
rect 14250 -4760 14370 -4720
rect 5960 -5404 6140 -5400
rect 5960 -5556 5974 -5404
rect 6126 -5556 6140 -5404
rect 5960 -5560 6140 -5556
rect 12020 -6440 12160 -6434
rect 11841 -6810 11850 -6730
rect 11930 -6810 11939 -6730
rect 7840 -7360 8240 -7340
rect 5144 -7490 5150 -7430
rect 5210 -7490 5216 -7430
rect 5334 -7434 5386 -7428
rect 5334 -7492 5386 -7486
rect 7840 -7500 7860 -7360
rect 8220 -7500 8240 -7360
rect 7840 -7520 8240 -7500
rect 11580 -7375 11770 -7360
rect 11580 -7525 11600 -7375
rect 11750 -7525 11770 -7375
rect 11580 -7540 11770 -7525
rect 9250 -7600 9350 -7580
rect 10010 -7600 10150 -7591
rect 8760 -7620 8820 -7614
rect 9250 -7620 9260 -7600
rect 8751 -7680 8760 -7620
rect 8820 -7670 9260 -7620
rect 9340 -7670 9350 -7600
rect 10000 -7660 10010 -7600
rect 8820 -7680 9350 -7670
rect 9450 -7670 10010 -7660
rect 8760 -7686 8820 -7680
rect 9450 -7730 9460 -7670
rect 9530 -7730 10010 -7670
rect 9450 -7740 10010 -7730
rect 11850 -7660 11930 -6810
rect 10150 -7740 11930 -7660
rect 10010 -7749 10150 -7740
rect 4135 -7780 9980 -7775
rect 10180 -7780 11695 -7775
rect 4135 -7885 11695 -7780
rect 11805 -7885 11811 -7775
rect 12020 -7970 12160 -6580
rect 15675 -6625 16025 -6515
rect 16135 -6625 16141 -6515
rect 15675 -7275 15785 -6625
rect 12275 -7385 15785 -7275
rect 12275 -7775 12385 -7385
rect 12275 -7891 12385 -7885
rect 3850 -8110 12160 -7970
rect 1880 -12030 14080 -11970
rect 1780 -12130 13090 -12070
rect 1680 -12230 12090 -12170
rect 1580 -12330 11090 -12270
rect 1480 -12430 10090 -12370
rect 1370 -12530 9090 -12470
rect 1270 -12630 8090 -12570
rect 1150 -12730 7090 -12670
rect 1030 -12830 6090 -12770
rect 930 -12930 4090 -12870
rect 810 -13030 3090 -12970
rect 690 -13130 2090 -13070
rect 590 -13230 1090 -13170
rect 1030 -13660 1090 -13230
rect 2030 -13660 2090 -13130
rect -10992 -13700 -10864 -13680
rect -10000 -13700 -9880 -13660
rect -9000 -13700 -8880 -13660
rect -8000 -13700 -7880 -13660
rect -7000 -13700 -6880 -13660
rect -6000 -13700 -5880 -13660
rect -5000 -13700 -4880 -13660
rect -4000 -13670 -3910 -13660
rect -4000 -13700 -3880 -13670
rect -3000 -13700 -2880 -13660
rect -2000 -13700 -1880 -13660
rect -1000 -13700 -880 -13660
rect 0 -13700 120 -13660
rect 1000 -13700 1120 -13660
rect 2000 -13670 2090 -13660
rect 3030 -13670 3090 -13030
rect 4030 -13670 4090 -12930
rect 5030 -13470 5150 -13410
rect 5210 -13470 5216 -13410
rect 5030 -13670 5090 -13470
rect 6030 -13670 6090 -12830
rect 7030 -13670 7090 -12730
rect 8030 -13670 8090 -12630
rect 9030 -13670 9090 -12530
rect 10030 -13670 10090 -12430
rect 11030 -13670 11090 -12330
rect 12030 -13670 12090 -12230
rect 13030 -13670 13090 -12130
rect 14020 -13670 14080 -12030
rect 14454 -13174 14506 -13168
rect 14506 -13220 17060 -13180
rect 14454 -13232 14506 -13226
rect 2000 -13700 2120 -13670
rect 3000 -13700 3120 -13670
rect 4000 -13700 4120 -13670
rect 5000 -13700 5120 -13670
rect 6000 -13700 6120 -13670
rect 7000 -13700 7120 -13670
rect 8000 -13700 8120 -13670
rect 9000 -13700 9120 -13670
rect 10000 -13700 10120 -13670
rect 11000 -13700 11120 -13670
rect 12000 -13700 12120 -13670
rect 13000 -13700 13120 -13670
rect 14000 -13700 14120 -13670
rect 15000 -13700 15120 -13670
rect 16000 -13700 16120 -13670
rect 17020 -13700 17060 -13220
rect -11400 -15200 -10600 -13700
rect -10300 -15200 -9500 -13700
rect -9300 -15200 -8500 -13700
rect -8300 -15200 -7500 -13700
rect -7300 -15200 -6500 -13700
rect -6300 -15200 -5500 -13700
rect -5300 -15200 -4500 -13700
rect -4300 -15200 -3500 -13700
rect -3300 -15200 -2500 -13700
rect -2300 -15200 -1500 -13700
rect -1300 -15200 -500 -13700
rect -300 -15200 500 -13700
rect 700 -15200 1500 -13700
rect 1700 -15200 2500 -13700
rect 2700 -15200 3500 -13700
rect 3700 -15200 4500 -13700
rect 4700 -15200 5500 -13700
rect 5700 -15200 6500 -13700
rect 6700 -15200 7500 -13700
rect 7700 -15200 8500 -13700
rect 8700 -15200 9500 -13700
rect 9700 -15200 10500 -13700
rect 10700 -15200 11500 -13700
rect 11700 -15200 12500 -13700
rect 12700 -15200 13500 -13700
rect 13700 -15200 14500 -13700
rect 14700 -13820 15500 -13700
rect 14700 -13880 15030 -13820
rect 15090 -13880 15500 -13820
rect 14700 -15200 15500 -13880
rect 15700 -13820 16500 -13700
rect 15700 -13880 16030 -13820
rect 16090 -13880 16500 -13820
rect 15700 -15200 16500 -13880
rect 16700 -15200 17500 -13700
<< via2 >>
rect 36 7588 92 7644
rect -1564 7524 -1508 7580
rect 1636 7572 1692 7628
rect 3236 7572 3292 7628
rect 4820 7556 4876 7612
rect 6436 7572 6492 7628
rect 8020 7572 8076 7628
rect 9700 7460 9756 7516
rect -4780 7316 -4724 7372
rect -652 7316 -596 7372
rect -6364 7140 -6308 7196
rect -7964 6948 -7908 7004
rect -11500 1300 -10900 1900
rect -12500 -100 -11900 500
rect -11500 -5100 -10850 -4450
rect 5810 6186 5870 6190
rect 5810 6134 5814 6186
rect 5814 6134 5866 6186
rect 5866 6134 5870 6186
rect 5810 6130 5870 6134
rect 4530 5978 4590 5982
rect 4530 5926 4534 5978
rect 4534 5926 4586 5978
rect 4586 5926 4590 5978
rect 4530 5922 4590 5926
rect -5036 5860 -4980 5916
rect -10400 -13520 -10336 -13456
rect 3234 5738 3294 5742
rect 3234 5686 3238 5738
rect 3238 5686 3290 5738
rect 3290 5686 3294 5738
rect 3234 5682 3294 5686
rect -654 5594 -594 5600
rect -654 5542 -650 5594
rect -650 5542 -598 5594
rect -598 5542 -594 5594
rect -654 5538 -594 5542
rect 1922 5562 1982 5566
rect 1922 5510 1926 5562
rect 1926 5510 1978 5562
rect 1978 5510 1982 5562
rect 1922 5506 1982 5510
rect -1934 5482 -1874 5486
rect -1934 5430 -1930 5482
rect -1930 5430 -1878 5482
rect -1878 5430 -1874 5482
rect -1934 5426 -1874 5430
rect 642 5402 702 5406
rect 642 5350 646 5402
rect 646 5350 698 5402
rect 698 5350 702 5402
rect 642 5346 702 5350
rect 7106 5466 7166 5470
rect 7106 5414 7110 5466
rect 7110 5414 7162 5466
rect 7162 5414 7166 5466
rect 7106 5410 7166 5414
rect 8386 5466 8446 5470
rect 8386 5414 8390 5466
rect 8390 5414 8442 5466
rect 8442 5414 8446 5466
rect 8386 5410 8446 5414
rect 9698 5466 9758 5470
rect 9698 5414 9702 5466
rect 9702 5414 9754 5466
rect 9754 5414 9758 5466
rect 9698 5410 9758 5414
rect -4490 5190 -4430 5250
rect -3214 5306 -3154 5310
rect -3214 5254 -3210 5306
rect -3210 5254 -3158 5306
rect -3158 5254 -3154 5306
rect -3214 5250 -3154 5254
rect -5160 3680 -5100 3740
rect -5060 3540 -5000 3600
rect -4960 3400 -4900 3460
rect -4860 3270 -4800 3330
rect 2352 3322 2408 3378
rect -4760 3130 -4700 3190
rect 2212 3192 2268 3248
rect 2072 3072 2128 3128
rect 1922 2982 1978 3038
rect 1750 2830 1810 2890
rect -3580 1920 -3500 2000
rect -2540 2060 -2460 2140
rect -345 1875 -215 2005
rect -1660 260 -1580 340
rect -1320 300 -1240 380
rect 4159 1360 4240 1441
rect 5215 1355 5285 1425
rect 379 674 501 796
rect 7270 280 7350 360
rect -2885 75 -2795 165
rect 655 -50 735 30
rect 2515 25 2585 95
rect -90 -180 10 -80
rect -300 -1660 -220 -1580
rect 8870 580 9050 760
rect 8900 -3220 9000 -3120
rect 11105 -4265 11275 -4095
rect 14575 -4555 14645 -4485
rect 14275 -4720 14345 -4650
rect 11850 -6810 11930 -6730
rect 7860 -7500 8220 -7360
rect 11605 -7520 11745 -7380
rect 8760 -7680 8820 -7620
rect 10010 -7740 10150 -7600
<< metal3 >>
rect -12510 17295 -12504 17905
rect -11894 17295 -11888 17905
rect -12503 505 -11896 17295
rect -11505 12901 -11499 13499
rect -10901 12901 -10895 13499
rect -11499 12580 -10901 12901
rect -11500 1905 -10900 12580
rect 31 7644 97 7649
rect 31 7588 36 7644
rect 92 7588 97 7644
rect -1569 7580 -1503 7585
rect 31 7583 97 7588
rect 1631 7628 1697 7633
rect -1569 7524 -1564 7580
rect -1508 7524 -1503 7580
rect -1569 7519 -1503 7524
rect -4785 7374 -4719 7377
rect -4785 7372 -1874 7374
rect -4785 7316 -4780 7372
rect -4724 7316 -1874 7372
rect -4785 7314 -1874 7316
rect -4785 7311 -4719 7314
rect -6369 7198 -6303 7201
rect -6369 7196 -3154 7198
rect -6369 7140 -6364 7196
rect -6308 7140 -3154 7196
rect -6369 7138 -3154 7140
rect -6369 7135 -6303 7138
rect -7969 7006 -7903 7009
rect -7969 7004 -4430 7006
rect -7969 6948 -7964 7004
rect -7908 6948 -4430 7004
rect -7969 6946 -4430 6948
rect -7969 6943 -7903 6946
rect -5041 5920 -4975 5921
rect -9696 5916 -4975 5920
rect -9696 5860 -5036 5916
rect -4980 5860 -4975 5916
rect -9696 5856 -4975 5860
rect -11505 1900 -10895 1905
rect -11505 1300 -11500 1900
rect -10900 1300 -10895 1900
rect -11505 1295 -10895 1300
rect -12505 500 -11895 505
rect -12505 -100 -12500 500
rect -11900 -100 -11895 500
rect -12505 -105 -11895 -100
rect -11600 -4445 -10700 -4300
rect -11600 -5105 -11505 -4445
rect -10845 -5105 -10700 -4445
rect -11600 -5200 -10700 -5105
rect -10405 -13456 -10331 -13451
rect -9696 -13456 -9632 5856
rect -5041 5855 -4975 5856
rect -4490 5255 -4430 6946
rect -3214 5328 -3154 7138
rect -1934 5504 -1874 7314
rect -1952 5486 -1856 5504
rect -1952 5426 -1934 5486
rect -1874 5426 -1856 5486
rect -1952 5424 -1856 5426
rect -1939 5421 -1869 5424
rect -1566 5406 -1506 7519
rect -657 7372 -591 7377
rect -657 7316 -652 7372
rect -596 7316 -591 7372
rect -657 7311 -591 7316
rect -654 5616 -594 7311
rect -672 5600 -576 5616
rect -672 5538 -654 5600
rect -594 5538 -576 5600
rect -672 5520 -576 5538
rect 34 5566 94 7583
rect 1631 7572 1636 7628
rect 1692 7572 1697 7628
rect 1631 7567 1697 7572
rect 3231 7628 3297 7633
rect 3231 7572 3236 7628
rect 3292 7572 3297 7628
rect 6431 7628 6497 7633
rect 3231 7567 3297 7572
rect 4815 7612 4881 7617
rect 1634 5742 1694 7567
rect 3234 5982 3294 7567
rect 4815 7556 4820 7612
rect 4876 7556 4881 7612
rect 6431 7572 6436 7628
rect 6492 7572 6497 7628
rect 6431 7567 6497 7572
rect 8015 7630 8081 7633
rect 8015 7628 8446 7630
rect 8015 7572 8020 7628
rect 8076 7572 8446 7628
rect 8015 7570 8446 7572
rect 8015 7567 8081 7570
rect 4815 7551 4881 7556
rect 4818 6190 4878 7551
rect 6434 7070 6494 7567
rect 6434 7010 7166 7070
rect 5792 6190 5888 6208
rect 4818 6130 5810 6190
rect 5870 6130 5888 6190
rect 5792 6112 5888 6130
rect 4512 5982 4608 6000
rect 3234 5922 4530 5982
rect 4590 5922 4608 5982
rect 4512 5904 4608 5922
rect 3216 5742 3312 5760
rect 1634 5682 3234 5742
rect 3294 5682 3312 5742
rect 3216 5664 3312 5682
rect 1904 5566 2000 5584
rect 34 5506 1922 5566
rect 1982 5506 2000 5566
rect 1904 5488 2000 5506
rect 7106 5488 7166 7010
rect 8386 5488 8446 7570
rect 9695 7516 9761 7521
rect 9695 7460 9700 7516
rect 9756 7460 9761 7516
rect 9695 7455 9761 7460
rect 7088 5470 7184 5488
rect 637 5406 707 5411
rect -1566 5346 642 5406
rect 702 5346 707 5406
rect 7088 5410 7106 5470
rect 7166 5410 7184 5470
rect 7088 5392 7184 5410
rect 8368 5470 8464 5488
rect 9698 5475 9758 7455
rect 8368 5410 8386 5470
rect 8446 5410 8464 5470
rect 8368 5392 8464 5410
rect 9693 5470 9763 5475
rect 9693 5410 9698 5470
rect 9758 5410 9763 5470
rect 9693 5405 9763 5410
rect 637 5341 707 5346
rect -3232 5310 -3136 5328
rect -4495 5250 -4425 5255
rect -4495 5190 -4490 5250
rect -4430 5190 -4425 5250
rect -3232 5250 -3214 5310
rect -3154 5250 -3136 5310
rect -3232 5216 -3136 5250
rect -4495 5185 -4425 5190
rect -5165 3740 -5095 3745
rect -5165 3680 -5160 3740
rect -5100 3680 2410 3740
rect -5165 3675 -5095 3680
rect -5065 3600 -4995 3605
rect -5065 3540 -5060 3600
rect -5000 3540 2270 3600
rect -5065 3535 -4995 3540
rect -4965 3460 -4895 3465
rect -4965 3400 -4960 3460
rect -4900 3400 2130 3460
rect -4965 3395 -4895 3400
rect -4865 3330 -4795 3335
rect -4865 3270 -4860 3330
rect -4800 3270 1980 3330
rect -4865 3265 -4795 3270
rect -4765 3190 -4695 3195
rect -4770 3130 -4760 3190
rect -4700 3130 1810 3190
rect -4765 3125 -4695 3130
rect 1750 2895 1810 3130
rect 1920 3050 1980 3270
rect 2070 3133 2130 3400
rect 2210 3253 2270 3540
rect 2350 3383 2410 3680
rect 2347 3378 2413 3383
rect 2347 3322 2352 3378
rect 2408 3322 2413 3378
rect 2347 3317 2413 3322
rect 2207 3248 2273 3253
rect 2207 3192 2212 3248
rect 2268 3192 2273 3248
rect 2207 3187 2273 3192
rect 2067 3128 2133 3133
rect 2067 3072 2072 3128
rect 2128 3072 2133 3128
rect 2067 3067 2133 3072
rect 1910 3038 1990 3050
rect 1910 2982 1922 3038
rect 1978 2982 1990 3038
rect 1910 2970 1990 2982
rect 1745 2890 1815 2895
rect 1745 2830 1750 2890
rect 1810 2830 1815 2890
rect 1745 2825 1815 2830
rect -2560 2145 -2440 2160
rect -2560 2055 -2545 2145
rect -2455 2055 -2440 2145
rect -2560 2040 -2440 2055
rect -3600 2005 -3480 2020
rect -3600 1915 -3585 2005
rect -3495 1915 -3480 2005
rect -3600 1900 -3480 1915
rect -380 2009 -180 2040
rect -380 1871 -349 2009
rect -211 1871 -180 2009
rect -380 1840 -180 1871
rect 4140 1445 4260 1460
rect 4140 1356 4155 1445
rect 4244 1356 4260 1445
rect 4140 1340 4260 1356
rect 5190 1429 5310 1450
rect 5190 1351 5211 1429
rect 5289 1351 5310 1429
rect 5190 1330 5310 1351
rect 374 796 396 801
rect 374 674 379 796
rect 374 669 396 674
rect 506 669 512 801
rect 8850 760 9070 780
rect 8850 580 8870 760
rect 9050 580 9070 760
rect 8850 560 9070 580
rect -1340 385 -1220 400
rect -1680 345 -1560 360
rect -1680 255 -1665 345
rect -1575 255 -1560 345
rect -1340 305 -1325 385
rect -1235 305 -1220 385
rect -1340 300 -1320 305
rect -1240 300 -1220 305
rect -1340 280 -1220 300
rect 7240 364 7370 380
rect 7240 276 7266 364
rect 7354 276 7370 364
rect 7240 260 7370 276
rect -1680 240 -1560 255
rect -2890 165 -2790 170
rect -2890 75 -2885 165
rect -2795 75 -2790 165
rect -2890 10 -2790 75
rect 2500 100 2600 110
rect 640 34 750 50
rect -2890 -75 10 10
rect 640 -54 651 34
rect 739 -54 750 34
rect 2500 20 2510 100
rect 2590 20 2600 100
rect 2500 10 2600 20
rect 640 -60 750 -54
rect -2890 -80 15 -75
rect -2890 -90 -90 -80
rect -95 -180 -90 -90
rect 10 -180 15 -80
rect -95 -185 15 -180
rect -392 -1560 -234 -1518
rect -392 -1575 -200 -1560
rect -392 -1665 -305 -1575
rect -215 -1665 -200 -1575
rect -392 -1680 -200 -1665
rect -392 -1686 -234 -1680
rect 8870 -3120 9050 560
rect 8870 -3220 8900 -3120
rect 9000 -3220 9050 -3120
rect 8870 -4090 9050 -3220
rect 11080 -4090 11300 -4070
rect 8870 -4095 11300 -4090
rect 8870 -4265 11105 -4095
rect 11275 -4265 11300 -4095
rect 8870 -4270 11300 -4265
rect 11080 -4290 11300 -4270
rect 13750 -4485 14650 -4480
rect 13750 -4555 14575 -4485
rect 14645 -4555 14650 -4485
rect 13750 -4560 14650 -4555
rect 13750 -4590 13830 -4560
rect 12210 -4670 13830 -4590
rect 14250 -4650 14370 -4630
rect 14250 -4655 14275 -4650
rect 14345 -4655 14370 -4650
rect 11845 -6730 11935 -6725
rect 12210 -6730 12290 -4670
rect 14250 -4725 14270 -4655
rect 14350 -4725 14370 -4655
rect 14250 -4760 14370 -4725
rect 11845 -6810 11850 -6730
rect 11930 -6810 12290 -6730
rect 11845 -6815 11935 -6810
rect 7840 -7360 8240 -7340
rect 7840 -7500 7860 -7360
rect 8220 -7500 8240 -7360
rect 7840 -7520 8240 -7500
rect 11580 -7376 11770 -7360
rect 11580 -7524 11601 -7376
rect 11749 -7524 11770 -7376
rect 11580 -7540 11770 -7524
rect 9980 -7595 10170 -7570
rect 8740 -7615 8840 -7600
rect 8740 -7685 8755 -7615
rect 8825 -7685 8840 -7615
rect 8740 -7700 8840 -7685
rect 9980 -7745 10005 -7595
rect 10155 -7745 10170 -7595
rect 9980 -7760 10170 -7745
rect -10405 -13520 -10400 -13456
rect -10336 -13520 -9632 -13456
rect -10405 -13525 -10331 -13520
<< via3 >>
rect -12504 17295 -11894 17905
rect -11499 12901 -10901 13499
rect -11505 -4450 -10845 -4445
rect -11505 -5100 -11500 -4450
rect -11500 -5100 -10850 -4450
rect -10850 -5100 -10845 -4450
rect -11505 -5105 -10845 -5100
rect -2545 2140 -2455 2145
rect -2545 2060 -2540 2140
rect -2540 2060 -2460 2140
rect -2460 2060 -2455 2140
rect -2545 2055 -2455 2060
rect -3585 2000 -3495 2005
rect -3585 1920 -3580 2000
rect -3580 1920 -3500 2000
rect -3500 1920 -3495 2000
rect -3585 1915 -3495 1920
rect -349 2005 -211 2009
rect -349 1875 -345 2005
rect -345 1875 -215 2005
rect -215 1875 -211 2005
rect -349 1871 -211 1875
rect 4155 1441 4244 1445
rect 4155 1360 4159 1441
rect 4159 1360 4240 1441
rect 4240 1360 4244 1441
rect 4155 1356 4244 1360
rect 5211 1425 5289 1429
rect 5211 1355 5215 1425
rect 5215 1355 5285 1425
rect 5285 1355 5289 1425
rect 5211 1351 5289 1355
rect 396 796 506 801
rect 396 674 501 796
rect 501 674 506 796
rect 396 669 506 674
rect -1665 340 -1575 345
rect -1665 260 -1660 340
rect -1660 260 -1580 340
rect -1580 260 -1575 340
rect -1665 255 -1575 260
rect -1325 380 -1235 385
rect -1325 305 -1320 380
rect -1320 305 -1240 380
rect -1240 305 -1235 380
rect 7266 360 7354 364
rect 7266 280 7270 360
rect 7270 280 7350 360
rect 7350 280 7354 360
rect 7266 276 7354 280
rect 651 30 739 34
rect 651 -50 655 30
rect 655 -50 735 30
rect 735 -50 739 30
rect 651 -54 739 -50
rect 2510 95 2590 100
rect 2510 25 2515 95
rect 2515 25 2585 95
rect 2585 25 2590 95
rect 2510 20 2590 25
rect -305 -1580 -215 -1575
rect -305 -1660 -300 -1580
rect -300 -1660 -220 -1580
rect -220 -1660 -215 -1580
rect -305 -1665 -215 -1660
rect 14270 -4720 14275 -4655
rect 14275 -4720 14345 -4655
rect 14345 -4720 14350 -4655
rect 14270 -4725 14350 -4720
rect 7860 -7500 8220 -7360
rect 11601 -7380 11749 -7376
rect 11601 -7520 11605 -7380
rect 11605 -7520 11745 -7380
rect 11745 -7520 11749 -7380
rect 11601 -7524 11749 -7520
rect 8755 -7620 8825 -7615
rect 8755 -7680 8760 -7620
rect 8760 -7680 8820 -7620
rect 8820 -7680 8825 -7620
rect 8755 -7685 8825 -7680
rect 10005 -7600 10155 -7595
rect 10005 -7740 10010 -7600
rect 10010 -7740 10150 -7600
rect 10150 -7740 10155 -7600
rect 10005 -7745 10155 -7740
<< metal4 >>
rect -13012 18000 16588 18420
rect -13012 17905 16600 18000
rect -13012 17616 -12504 17905
rect -13000 17450 -12504 17616
rect -13012 17295 -12504 17450
rect -11894 17450 16600 17905
rect -11894 17295 16608 17450
rect -13012 16960 16608 17295
rect -11622 13544 17998 14034
rect -11600 13499 17988 13544
rect -11600 12901 -11499 13499
rect -10901 12901 17988 13499
rect -11600 12878 17988 12901
rect -11612 12388 18008 12878
rect -2546 2145 -2454 2146
rect -2546 2055 -2545 2145
rect -2455 2140 -2454 2145
rect -2455 2060 -1240 2140
rect -2455 2055 -2454 2060
rect -2546 2054 -2454 2055
rect -3586 2005 -3494 2006
rect -3586 1915 -3585 2005
rect -3495 2000 -3494 2005
rect -3495 1920 -2660 2000
rect -3495 1915 -3494 1920
rect -3586 1914 -3494 1915
rect -2740 1640 -2660 1920
rect -1320 1740 -1240 2060
rect 384 2124 2635 2215
rect -350 2009 -120 2010
rect -350 1871 -349 2009
rect -211 2008 -120 2009
rect 384 2008 475 2124
rect -211 1917 475 2008
rect -211 1910 -120 1917
rect -211 1871 -210 1910
rect -1660 346 -1580 800
rect -1320 386 -1240 600
rect -1326 385 -1234 386
rect -1666 345 -1574 346
rect -1666 255 -1665 345
rect -1575 255 -1574 345
rect -1326 305 -1325 385
rect -1235 305 -1234 385
rect -1326 304 -1234 305
rect -1666 254 -1574 255
rect -350 -1420 -210 1871
rect 2544 1446 2635 2124
rect 2544 1445 4245 1446
rect 2544 1356 4155 1445
rect 4244 1356 4245 1445
rect 5190 1430 5310 1450
rect 2544 1355 4245 1356
rect 4380 1429 5310 1430
rect 4380 1351 5211 1429
rect 5289 1351 5310 1429
rect 4380 1350 5310 1351
rect 4380 1270 4460 1350
rect 5190 1330 5310 1350
rect 2510 1190 4460 1270
rect 395 801 507 802
rect 395 669 396 801
rect 506 790 507 801
rect 506 680 1015 790
rect 506 669 507 680
rect 395 668 507 669
rect 650 34 740 210
rect 2510 101 2590 1190
rect 7265 364 8585 365
rect 7265 276 7266 364
rect 7354 276 8585 364
rect 7265 275 8585 276
rect 650 -54 651 34
rect 739 -54 740 34
rect 2509 100 2591 101
rect 2509 20 2510 100
rect 2590 20 2591 100
rect 2509 19 2591 20
rect 650 -55 740 -54
rect 2514 -804 2586 19
rect 2514 -876 4026 -804
rect 3954 -1136 4026 -876
rect -360 -1520 -200 -1420
rect -560 -1575 -200 -1520
rect -560 -1665 -305 -1575
rect -215 -1665 -200 -1575
rect -560 -1700 -200 -1665
rect 8495 -2405 8585 275
rect 8420 -2495 8585 -2405
rect -11600 -4445 -10700 -4300
rect -11600 -5105 -11505 -4445
rect -10845 -5105 -10700 -4445
rect -11600 -5200 -10700 -5105
rect -11500 -5725 -10845 -5200
rect -11500 -13600 -10880 -5725
rect 8420 -6230 8510 -2495
rect 14269 -4655 14351 -4654
rect 14269 -4725 14270 -4655
rect 14350 -4725 14351 -4655
rect 14269 -4726 14351 -4725
rect 14275 -5525 14345 -4726
rect 12815 -5595 14345 -5525
rect 12815 -5815 12885 -5595
rect 8420 -6240 8570 -6230
rect 8420 -6380 8820 -6240
rect 8420 -6480 8540 -6380
rect 8420 -7340 8520 -6480
rect 7840 -7360 8240 -7340
rect 7840 -7500 7860 -7360
rect 8220 -7500 8240 -7360
rect 7840 -7520 8240 -7500
rect 7840 -7940 7940 -7520
rect 8400 -7620 8520 -7340
rect 11580 -7376 11770 -7360
rect 11580 -7524 11601 -7376
rect 11749 -7524 11770 -7376
rect 11580 -7540 11770 -7524
rect 9980 -7595 10170 -7570
rect 8754 -7615 8826 -7614
rect 8754 -7620 8755 -7615
rect 8400 -7680 8755 -7620
rect 8754 -7685 8755 -7680
rect 8825 -7685 8826 -7615
rect 8754 -7686 8826 -7685
rect 9980 -7745 10005 -7595
rect 10155 -7745 10170 -7595
rect 9980 -7760 10170 -7745
rect 10010 -8920 10150 -7760
rect 11600 -8750 11690 -7540
rect -11900 -14584 -7400 -13600
rect -11906 -14600 -7400 -14584
rect -11906 -15098 -7406 -14600
use sky130_fd_pr__cap_mim_m3_1_VT6YF8  C1
timestamp 1667918091
transform 1 0 -2070 0 1 1200
box -850 -700 849 700
use sky130_fd_pr__cap_mim_m3_1_AFDLP7  C2
timestamp 1667918091
transform 0 1 1520 -1 0 1079
box -950 -900 949 900
use sky130_fd_pr__cap_mim_m3_1_AFDLP7  C3
timestamp 1667918091
transform 1 0 10740 0 1 -9520
box -950 -900 949 900
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  C4
timestamp 1667918091
transform 1 0 6350 0 1 -9700
box -2150 -2100 2149 2100
use CurrentMirror_post  CurrentMirror_post_0
timestamp 1667225002
transform 1 0 -4260 0 1 -6200
box 460 480 8480 1932
use CurrentMirror_post  CurrentMirror_post_1
timestamp 1667225002
transform 1 0 -4260 0 1 -7680
box 460 480 8480 1932
use Inverter_post  Inverter_post_0
timestamp 1667917589
transform 1 0 12564 0 1 -4190
box -624 -240 -128 896
use Inverter_post  Inverter_post_1
timestamp 1667917589
transform -1 0 8882 0 1 1810
box -624 -240 -128 896
use sky130_fd_pr__nfet_01v8_lvt_KP8PNM  M6
timestamp 1667938751
transform 1 0 6026 0 1 -6801
box -1586 -399 1586 399
use sky130_fd_pr__nfet_01v8_lvt_MHJ2VF  M7
timestamp 1667938751
transform 1 0 7896 0 1 -6921
box -296 -279 296 279
use sky130_fd_pr__pfet_01v8_lvt_8MQB6L  M8
timestamp 1667938215
transform -1 0 6026 0 -1 -5996
box -1586 -404 1586 404
use sky130_fd_pr__pfet_01v8_lvt_7PDTEF  M9
timestamp 1667938215
transform -1 0 7896 0 -1 -6116
box -296 -284 296 284
use M  M_0
timestamp 1667919441
transform 1 0 -227 0 1 2453
box -53 -53 517 505
use M  M_1
timestamp 1667919441
transform -1 0 797 0 -1 2905
box -53 -53 517 505
use M  M_3
timestamp 1667919441
transform -1 0 517 0 -1 -1415
box -53 -53 517 505
use M  M_4
timestamp 1667919441
transform -1 0 9727 0 -1 -7235
box -53 -53 517 505
use M  M_5
timestamp 1667919441
transform -1 0 9157 0 -1 -7235
box -53 -53 517 505
use M  M_11
timestamp 1667919441
transform 0 -1 -4435 1 0 4793
box -53 -53 517 505
use OTA_post  OTA_post_0
timestamp 1668277347
transform 1 0 -4560 0 1 -3320
box 560 820 4240 3330
use OTA_post  OTA_post_1
timestamp 1668277347
transform 1 0 140 0 1 -3320
box 560 820 4240 3330
use OTA_post  OTA_post_2
timestamp 1668277347
transform 1 0 4190 0 1 -3320
box 560 820 4240 3330
use OTA_post  OTA_post_3
timestamp 1668277347
transform -1 0 12720 0 1 -8020
box 560 820 4240 3330
use OTA_post  OTA_post_4
timestamp 1668277347
transform -1 0 16690 0 1 -8020
box 560 820 4240 3330
use Tgate_post  Tgate_post_0
timestamp 1667228915
transform 1 0 -1900 0 1 240
box -1080 420 -10 1600
use Tgate_post  Tgate_post_1
timestamp 1667228915
transform 1 0 -2940 0 1 240
box -1080 420 -10 1600
use Tgate_post  Tgate_post_2
timestamp 1667228915
transform 1 0 -860 0 1 240
box -1080 420 -10 1600
use Tgate_post  Tgate_post_3
timestamp 1667228915
transform 1 0 180 0 1 240
box -1080 420 -10 1600
use Tgate_post  Tgate_post_4
timestamp 1667228915
transform 1 0 8990 0 1 1130
box -1080 420 -10 1600
use Tgate_post  Tgate_post_5
timestamp 1667228915
transform 1 0 4800 0 1 1130
box -1080 420 -10 1600
use Tgate_post  Tgate_post_6
timestamp 1667228915
transform 1 0 5850 0 1 1130
box -1080 420 -10 1600
use Tgate_post  Tgate_post_7
timestamp 1667228915
transform 1 0 7940 0 1 1130
box -1080 420 -10 1600
use Tgate_post  Tgate_post_8
timestamp 1667228915
transform 1 0 6900 0 1 1130
box -1080 420 -10 1600
use Tgate_post  Tgate_post_10
timestamp 1667228915
transform 1 0 13530 0 1 -4870
box -1080 420 -10 1600
use Tgate_post  Tgate_post_11
timestamp 1667228915
transform 1 0 14580 0 1 -4870
box -1080 420 -10 1600
use VoltageDivider-P_post  VoltageDivider-P_post_0
timestamp 1667915364
transform 1 0 7580 0 1 -5050
box -980 -300 512 1128
<< labels >>
flabel via2 -11500 1500 -11500 1500 0 FreeSans 1600 0 0 0 VDD
port 1 nsew power input
flabel metal2 5060 -14460 5060 -14460 0 FreeSans 1600 90 0 0 Vref_sel_c
port 54 nsew signal input
flabel metal2 -11460 -6060 -11460 -6060 0 FreeSans 1600 0 0 0 pd12_b
port 53 nsew signal input
flabel metal2 -11460 -7060 -11460 -7060 0 FreeSans 1600 0 0 0 pd12_a
port 52 nsew signal input
flabel metal2 9660 8480 9660 8480 0 FreeSans 1600 0 0 0 PD12
port 51 nsew signal output
flabel metal2 -11460 -8060 -11460 -8060 0 FreeSans 1600 0 0 0 pd11_b
port 50 nsew signal input
flabel metal2 -11460 -9060 -11460 -9060 0 FreeSans 1600 0 0 0 pd11_a
port 49 nsew signal input
flabel metal2 8060 8480 8060 8480 0 FreeSans 1600 0 0 0 PD11
port 48 nsew signal output
flabel metal2 -11440 -10060 -11440 -10060 0 FreeSans 1600 0 0 0 pd10_b
port 47 nsew signal input
flabel metal2 -11460 -11060 -11460 -11060 0 FreeSans 1600 0 0 0 pd10_a
port 46 nsew signal input
flabel metal2 6460 8480 6460 8480 0 FreeSans 1600 0 0 0 PD10
port 45 nsew signal output
flabel metal2 -11440 -12060 -11440 -12060 0 FreeSans 1600 0 0 0 pd9_b
port 44 nsew signal input
flabel metal2 -11460 -13060 -11460 -13060 0 FreeSans 1600 0 0 0 pd9_a
port 43 nsew signal input
flabel metal2 4860 8480 4860 8480 0 FreeSans 1600 0 0 0 PD9
port 42 nsew signal output
flabel metal2 -10940 -14460 -10940 -14460 0 FreeSans 1600 90 0 0 pd8_b
port 41 nsew signal input
flabel metal2 -9940 -14460 -9940 -14460 0 FreeSans 1600 90 0 0 pd8_a
port 40 nsew signal input
flabel metal2 3260 8480 3260 8480 0 FreeSans 1600 0 0 0 PD8
port 39 nsew signal output
flabel metal2 -8940 -14460 -8940 -14460 0 FreeSans 1600 90 0 0 pd7_b
port 38 nsew signal input
flabel metal2 -7940 -14460 -7940 -14460 0 FreeSans 1600 90 0 0 pd7_a
port 37 nsew signal input
flabel metal2 1660 8480 1660 8480 0 FreeSans 1600 0 0 0 PD7
port 35 nsew signal output
flabel metal2 -6940 -14460 -6940 -14460 0 FreeSans 1600 90 0 0 pd6_b
port 34 nsew signal input
flabel metal2 -5940 -14460 -5940 -14460 0 FreeSans 1600 90 0 0 pd6_a
port 33 nsew signal input
flabel metal2 60 8480 60 8480 0 FreeSans 1600 0 0 0 PD6
port 32 nsew signal output
flabel metal2 -4940 -14460 -4940 -14460 0 FreeSans 1600 90 0 0 pd5_b
port 31 nsew signal input
flabel metal2 -3940 -14460 -3940 -14460 0 FreeSans 1600 90 0 0 pd5_a
port 30 nsew signal input
flabel metal2 -1540 8480 -1540 8480 0 FreeSans 1600 0 0 0 PD5
port 29 nsew signal output
flabel metal2 -2940 -14460 -2940 -14460 0 FreeSans 1600 90 0 0 pd4_b
port 28 nsew signal input
flabel metal2 -1940 -14460 -1940 -14460 0 FreeSans 1600 90 0 0 pd4_a
port 27 nsew signal input
flabel metal2 -3140 8480 -3140 8480 0 FreeSans 1600 0 0 0 PD4
port 26 nsew signal output
flabel metal2 -940 -14460 -940 -14460 0 FreeSans 1600 90 0 0 pd3_b
port 25 nsew signal input
flabel metal2 60 -14460 60 -14460 0 FreeSans 1600 90 0 0 pd3_a
port 24 nsew signal input
flabel metal2 -4740 8480 -4740 8480 0 FreeSans 1600 0 0 0 PD3
port 23 nsew signal output
flabel metal2 1060 -14460 1060 -14460 0 FreeSans 1600 90 0 0 pd2_b
port 22 nsew signal input
flabel metal2 2060 -14460 2060 -14460 0 FreeSans 1600 90 0 0 pd2_a
port 21 nsew signal input
flabel metal2 -6340 8480 -6340 8480 0 FreeSans 1600 0 0 0 PD2
port 20 nsew signal output
flabel metal2 10060 -14460 10060 -14460 0 FreeSans 1600 90 0 0 CMP_out_c
port 19 nsew signal input
flabel metal2 9060 -14460 9060 -14460 0 FreeSans 1600 90 0 0 OTA_sh_c
port 18 nsew signal input
flabel metal2 8060 -14460 8060 -14460 0 FreeSans 1600 90 0 0 Vref_cmp_c
port 17 nsew signal input
flabel metal2 7060 -14460 7060 -14460 0 FreeSans 1600 90 0 0 SH_out_c
port 16 nsew signal input
flabel metal2 6060 -14460 6060 -14460 0 FreeSans 1600 90 0 0 OTA_out_c
port 15 nsew signal input
flabel metal2 15060 -14440 15060 -14440 0 FreeSans 1600 90 0 0 sh_rst
port 14 nsew signal input
flabel metal2 16060 -14460 16060 -14460 0 FreeSans 1600 90 0 0 sh_cmp
port 13 nsew signal input
flabel metal2 17060 -14460 17060 -14460 0 FreeSans 1600 90 0 0 sh
port 12 nsew signal input
flabel metal2 13060 -14460 13060 -14460 0 FreeSans 1600 0 0 0 sw2
port 10 nsew signal input
flabel metal2 14060 -14460 14060 -14460 0 FreeSans 1600 0 0 0 sw1
port 9 nsew signal input
flabel metal2 12060 -14460 12060 -14460 0 FreeSans 1600 0 0 0 Vd2
port 8 nsew signal input
flabel metal2 11060 -14460 11060 -14460 0 FreeSans 1600 0 0 0 Vd1
port 7 nsew signal input
flabel via2 -11480 -4640 -11480 -4640 0 FreeSans 1600 0 0 0 Ibias
port 6 nsew power input
flabel metal2 3060 -14460 3060 -14460 0 FreeSans 1600 0 0 0 pd1_b
port 5 nsew signal input
flabel metal2 4060 -14460 4060 -14460 0 FreeSans 1600 0 0 0 pd1_a
port 4 nsew signal input
flabel metal2 -7940 8480 -7940 8480 0 FreeSans 1600 0 0 0 PD1
port 3 nsew signal output
flabel metal2 -11500 200 -11500 200 0 FreeSans 1600 0 0 0 VSS
port 2 nsew ground input
flabel metal2 16500 1360 16500 1360 0 FreeSans 1600 0 0 0 Aout
port 0 nsew signal output
flabel metal2 16400 0 16400 0 0 FreeSans 1600 0 0 0 CMP
port 55 nsew signal output
<< end >>
