magic
tech sky130A
magscale 1 2
timestamp 1678372745
<< dnwell >>
rect 30500 5100 49800 6500
rect 30500 1900 37500 5100
rect 42700 1900 49800 5100
rect 30500 500 49800 1900
rect 60500 5100 79800 6500
rect 60500 1900 67500 5100
rect 72700 1900 79800 5100
rect 60500 500 79800 1900
rect 90500 5100 109800 6500
rect 90500 1900 97500 5100
rect 102700 1900 109800 5100
rect 90500 500 109800 1900
rect 120500 5100 139800 6500
rect 120500 1900 127500 5100
rect 132700 1900 139800 5100
rect 120500 500 139800 1900
rect 150500 5100 169800 6500
rect 150500 1900 157500 5100
rect 162700 1900 169800 5100
rect 150500 500 169800 1900
rect 180500 5100 199800 6500
rect 180500 1900 187500 5100
rect 192700 1900 199800 5100
rect 180500 500 199800 1900
rect 210500 5100 229800 6500
rect 210500 1900 217500 5100
rect 222700 1900 229800 5100
rect 210500 500 229800 1900
rect 240500 5100 259800 6500
rect 240500 1900 247500 5100
rect 252700 1900 259800 5100
rect 240500 500 259800 1900
rect 270500 5100 289800 6500
rect 270500 1900 277500 5100
rect 282700 1900 289800 5100
rect 270500 500 289800 1900
rect 300500 5100 319800 6500
rect 300500 1900 307500 5100
rect 312700 1900 319800 5100
rect 300500 500 319800 1900
rect 330500 5100 349800 6500
rect 330500 1900 337500 5100
rect 342700 1900 349800 5100
rect 330500 500 349800 1900
rect 360500 5100 379800 6500
rect 360500 1900 367500 5100
rect 372700 1900 379800 5100
rect 360500 500 379800 1900
<< photodiode >>
rect 39700 3300 40300 3900
rect 69700 3300 70300 3900
rect 99700 3300 100300 3900
rect 129700 3300 130300 3900
rect 159700 3300 160300 3900
rect 189700 3300 190300 3900
rect 219700 3300 220300 3900
rect 249700 3300 250300 3900
rect 279700 3300 280300 3900
rect 309700 3300 310300 3900
rect 339700 3300 340300 3900
rect 369700 3300 370300 3900
<< nwell >>
rect 30300 6100 50000 6700
rect 30300 900 30900 6100
rect 37100 5000 43100 5500
rect 37100 2000 37600 5000
rect 39860 3460 40140 3740
rect 42600 2000 43100 5000
rect 37100 1500 43100 2000
rect 49400 900 50000 6100
rect 30300 300 50000 900
rect 60300 6100 80000 6700
rect 60300 900 60900 6100
rect 67100 5000 73100 5500
rect 67100 2000 67600 5000
rect 69860 3460 70140 3740
rect 72600 2000 73100 5000
rect 67100 1500 73100 2000
rect 79400 900 80000 6100
rect 60300 300 80000 900
rect 90300 6100 110000 6700
rect 90300 900 91500 6100
rect 97100 5000 103100 5500
rect 97100 2000 97600 5000
rect 99860 3460 100140 3740
rect 102600 2000 103100 5000
rect 97100 1500 103100 2000
rect 108800 900 110000 6100
rect 90300 300 110000 900
rect 120300 6100 140000 6700
rect 120300 900 121500 6100
rect 127100 5000 133100 5500
rect 127100 2000 127600 5000
rect 129860 3460 130140 3740
rect 132600 2000 133100 5000
rect 127100 1500 133100 2000
rect 138800 900 140000 6100
rect 120300 300 140000 900
rect 150300 6100 170000 6700
rect 150300 900 152100 6100
rect 157100 5000 163100 5500
rect 157100 2000 157600 5000
rect 159860 3460 160140 3740
rect 162600 2000 163100 5000
rect 157100 1500 163100 2000
rect 168200 900 170000 6100
rect 150300 300 170000 900
rect 180300 6100 200000 6700
rect 180300 900 182100 6100
rect 187100 5000 193100 5500
rect 187100 2000 187600 5000
rect 189860 3460 190140 3740
rect 192600 2000 193100 5000
rect 187100 1500 193100 2000
rect 198200 900 200000 6100
rect 180300 300 200000 900
rect 210300 6100 230000 6700
rect 210300 900 212700 6100
rect 217100 5000 223100 5500
rect 217100 2000 217600 5000
rect 219860 3460 220140 3740
rect 222600 2000 223100 5000
rect 217100 1500 223100 2000
rect 227600 900 230000 6100
rect 210300 300 230000 900
rect 240300 6100 260000 6700
rect 240300 900 242700 6100
rect 247100 5000 253100 5500
rect 247100 2000 247600 5000
rect 249860 3460 250140 3740
rect 252600 2000 253100 5000
rect 247100 1500 253100 2000
rect 257600 900 260000 6100
rect 240300 300 260000 900
rect 270300 6100 290000 6700
rect 270300 900 273300 6100
rect 277100 5000 283100 5500
rect 277100 2000 277600 5000
rect 279860 3460 280140 3740
rect 282600 2000 283100 5000
rect 277100 1500 283100 2000
rect 287000 900 290000 6100
rect 270300 300 290000 900
rect 300300 6100 320000 6700
rect 300300 900 303300 6100
rect 307100 5000 313100 5500
rect 307100 2000 307600 5000
rect 309860 3460 310140 3740
rect 312600 2000 313100 5000
rect 307100 1500 313100 2000
rect 317000 900 320000 6100
rect 300300 300 320000 900
rect 330300 6100 350000 6700
rect 330300 900 333900 6100
rect 337100 5000 343100 5500
rect 337100 2000 337600 5000
rect 339860 3460 340140 3740
rect 342600 2000 343100 5000
rect 337100 1500 343100 2000
rect 346400 900 350000 6100
rect 330300 300 350000 900
rect 360300 6100 380000 6700
rect 360300 900 363900 6100
rect 367100 5000 373100 5500
rect 367100 2000 367600 5000
rect 369860 3460 370140 3740
rect 372600 2000 373100 5000
rect 367100 1500 373100 2000
rect 376400 900 380000 6100
rect 360300 300 380000 900
<< pwell >>
rect 30000 6700 50300 7000
rect 30000 300 30300 6700
rect 50000 300 50300 6700
rect 30000 0 50300 300
rect 60000 6700 80300 7000
rect 60000 300 60300 6700
rect 80000 300 80300 6700
rect 60000 0 80300 300
rect 90000 6700 110300 7000
rect 90000 300 90300 6700
rect 110000 300 110300 6700
rect 90000 0 110300 300
rect 120000 6700 140300 7000
rect 120000 300 120300 6700
rect 140000 300 140300 6700
rect 120000 0 140300 300
rect 150000 6700 170300 7000
rect 150000 300 150300 6700
rect 170000 300 170300 6700
rect 150000 0 170300 300
rect 180000 6700 200300 7000
rect 180000 300 180300 6700
rect 200000 300 200300 6700
rect 180000 0 200300 300
rect 210000 6700 230300 7000
rect 210000 300 210300 6700
rect 230000 300 230300 6700
rect 210000 0 230300 300
rect 240000 6700 260300 7000
rect 240000 300 240300 6700
rect 260000 300 260300 6700
rect 240000 0 260300 300
rect 270000 6700 290300 7000
rect 270000 300 270300 6700
rect 290000 300 290300 6700
rect 270000 0 290300 300
rect 300000 6700 320300 7000
rect 300000 300 300300 6700
rect 320000 300 320300 6700
rect 300000 0 320300 300
rect 330000 6700 350300 7000
rect 330000 300 330300 6700
rect 350000 300 350300 6700
rect 330000 0 350300 300
rect 360000 6700 380300 7000
rect 360000 300 360300 6700
rect 380000 300 380300 6700
rect 360000 0 380300 300
<< psubdiff >>
rect 30100 6800 30300 6900
rect 50000 6800 50200 6900
rect 30100 6700 30200 6800
rect 50100 6700 50200 6800
rect 30100 200 30200 300
rect 50100 200 50200 300
rect 30100 100 30300 200
rect 50000 100 50200 200
rect 60100 6800 60300 6900
rect 80000 6800 80200 6900
rect 60100 6700 60200 6800
rect 80100 6700 80200 6800
rect 60100 200 60200 300
rect 80100 200 80200 300
rect 60100 100 60300 200
rect 80000 100 80200 200
rect 90100 6800 90300 6900
rect 110000 6800 110200 6900
rect 90100 6700 90200 6800
rect 110100 6700 110200 6800
rect 90100 200 90200 300
rect 110100 200 110200 300
rect 90100 100 90300 200
rect 110000 100 110200 200
rect 120100 6800 120300 6900
rect 140000 6800 140200 6900
rect 120100 6700 120200 6800
rect 140100 6700 140200 6800
rect 120100 200 120200 300
rect 140100 200 140200 300
rect 120100 100 120300 200
rect 140000 100 140200 200
rect 150100 6800 150300 6900
rect 170000 6800 170200 6900
rect 150100 6700 150200 6800
rect 170100 6700 170200 6800
rect 150100 200 150200 300
rect 170100 200 170200 300
rect 150100 100 150300 200
rect 170000 100 170200 200
rect 180100 6800 180300 6900
rect 200000 6800 200200 6900
rect 180100 6700 180200 6800
rect 200100 6700 200200 6800
rect 180100 200 180200 300
rect 200100 200 200200 300
rect 180100 100 180300 200
rect 200000 100 200200 200
rect 210100 6800 210300 6900
rect 230000 6800 230200 6900
rect 210100 6700 210200 6800
rect 230100 6700 230200 6800
rect 210100 200 210200 300
rect 230100 200 230200 300
rect 210100 100 210300 200
rect 230000 100 230200 200
rect 240100 6800 240300 6900
rect 260000 6800 260200 6900
rect 240100 6700 240200 6800
rect 260100 6700 260200 6800
rect 240100 200 240200 300
rect 260100 200 260200 300
rect 240100 100 240300 200
rect 260000 100 260200 200
rect 270100 6800 270300 6900
rect 290000 6800 290200 6900
rect 270100 6700 270200 6800
rect 290100 6700 290200 6800
rect 270100 200 270200 300
rect 290100 200 290200 300
rect 270100 100 270300 200
rect 290000 100 290200 200
rect 300100 6800 300300 6900
rect 320000 6800 320200 6900
rect 300100 6700 300200 6800
rect 320100 6700 320200 6800
rect 300100 200 300200 300
rect 320100 200 320200 300
rect 300100 100 300300 200
rect 320000 100 320200 200
rect 330100 6800 330300 6900
rect 350000 6800 350200 6900
rect 330100 6700 330200 6800
rect 350100 6700 350200 6800
rect 330100 200 330200 300
rect 350100 200 350200 300
rect 330100 100 330300 200
rect 350000 100 350200 200
rect 360100 6800 360300 6900
rect 380000 6800 380200 6900
rect 360100 6700 360200 6800
rect 380100 6700 380200 6800
rect 360100 200 360200 300
rect 380100 200 380200 300
rect 360100 100 360300 200
rect 380000 100 380200 200
<< nsubdiff >>
rect 30500 6300 30700 6500
rect 39300 6300 39500 6500
rect 40500 6300 40700 6500
rect 49600 6300 49800 6500
rect 37300 3900 37500 4300
rect 42700 3900 42900 4300
rect 39920 3640 40080 3680
rect 39920 3560 39960 3640
rect 40040 3560 40080 3640
rect 39920 3520 40080 3560
rect 37300 2900 37500 3300
rect 42700 2900 42900 3300
rect 30500 500 30700 700
rect 39300 500 39500 700
rect 40500 500 40700 700
rect 49600 500 49800 700
rect 60500 6300 60700 6500
rect 69300 6300 69500 6500
rect 70500 6300 70700 6500
rect 79600 6300 79800 6500
rect 67300 3900 67500 4300
rect 72700 3900 72900 4300
rect 69920 3640 70080 3680
rect 69920 3560 69960 3640
rect 70040 3560 70080 3640
rect 69920 3520 70080 3560
rect 67300 2900 67500 3300
rect 72700 2900 72900 3300
rect 60500 500 60700 700
rect 69300 500 69500 700
rect 70500 500 70700 700
rect 79600 500 79800 700
rect 90500 6300 90700 6500
rect 99300 6300 99500 6500
rect 100500 6300 100700 6500
rect 109600 6300 109800 6500
rect 97300 3900 97500 4300
rect 102700 3900 102900 4300
rect 99920 3640 100080 3680
rect 99920 3560 99960 3640
rect 100040 3560 100080 3640
rect 99920 3520 100080 3560
rect 97300 2900 97500 3300
rect 102700 2900 102900 3300
rect 90500 500 90700 700
rect 99300 500 99500 700
rect 100500 500 100700 700
rect 109600 500 109800 700
rect 120500 6300 120700 6500
rect 129300 6300 129500 6500
rect 130500 6300 130700 6500
rect 139600 6300 139800 6500
rect 127300 3900 127500 4300
rect 132700 3900 132900 4300
rect 129920 3640 130080 3680
rect 129920 3560 129960 3640
rect 130040 3560 130080 3640
rect 129920 3520 130080 3560
rect 127300 2900 127500 3300
rect 132700 2900 132900 3300
rect 120500 500 120700 700
rect 129300 500 129500 700
rect 130500 500 130700 700
rect 139600 500 139800 700
rect 150500 6300 150700 6500
rect 159300 6300 159500 6500
rect 160500 6300 160700 6500
rect 169600 6300 169800 6500
rect 157300 3900 157500 4300
rect 162700 3900 162900 4300
rect 159920 3640 160080 3680
rect 159920 3560 159960 3640
rect 160040 3560 160080 3640
rect 159920 3520 160080 3560
rect 157300 2900 157500 3300
rect 162700 2900 162900 3300
rect 150500 500 150700 700
rect 159300 500 159500 700
rect 160500 500 160700 700
rect 169600 500 169800 700
rect 180500 6300 180700 6500
rect 189300 6300 189500 6500
rect 190500 6300 190700 6500
rect 199600 6300 199800 6500
rect 187300 3900 187500 4300
rect 192700 3900 192900 4300
rect 189920 3640 190080 3680
rect 189920 3560 189960 3640
rect 190040 3560 190080 3640
rect 189920 3520 190080 3560
rect 187300 2900 187500 3300
rect 192700 2900 192900 3300
rect 180500 500 180700 700
rect 189300 500 189500 700
rect 190500 500 190700 700
rect 199600 500 199800 700
rect 210500 6300 210700 6500
rect 219300 6300 219500 6500
rect 220500 6300 220700 6500
rect 229600 6300 229800 6500
rect 217300 3900 217500 4300
rect 222700 3900 222900 4300
rect 219920 3640 220080 3680
rect 219920 3560 219960 3640
rect 220040 3560 220080 3640
rect 219920 3520 220080 3560
rect 217300 2900 217500 3300
rect 222700 2900 222900 3300
rect 210500 500 210700 700
rect 219300 500 219500 700
rect 220500 500 220700 700
rect 229600 500 229800 700
rect 240500 6300 240700 6500
rect 249300 6300 249500 6500
rect 250500 6300 250700 6500
rect 259600 6300 259800 6500
rect 247300 3900 247500 4300
rect 252700 3900 252900 4300
rect 249920 3640 250080 3680
rect 249920 3560 249960 3640
rect 250040 3560 250080 3640
rect 249920 3520 250080 3560
rect 247300 2900 247500 3300
rect 252700 2900 252900 3300
rect 240500 500 240700 700
rect 249300 500 249500 700
rect 250500 500 250700 700
rect 259600 500 259800 700
rect 270500 6300 270700 6500
rect 279300 6300 279500 6500
rect 280500 6300 280700 6500
rect 289600 6300 289800 6500
rect 277300 3900 277500 4300
rect 282700 3900 282900 4300
rect 279920 3640 280080 3680
rect 279920 3560 279960 3640
rect 280040 3560 280080 3640
rect 279920 3520 280080 3560
rect 277300 2900 277500 3300
rect 282700 2900 282900 3300
rect 270500 500 270700 700
rect 279300 500 279500 700
rect 280500 500 280700 700
rect 289600 500 289800 700
rect 300500 6300 300700 6500
rect 309300 6300 309500 6500
rect 310500 6300 310700 6500
rect 319600 6300 319800 6500
rect 307300 3900 307500 4300
rect 312700 3900 312900 4300
rect 309920 3640 310080 3680
rect 309920 3560 309960 3640
rect 310040 3560 310080 3640
rect 309920 3520 310080 3560
rect 307300 2900 307500 3300
rect 312700 2900 312900 3300
rect 300500 500 300700 700
rect 309300 500 309500 700
rect 310500 500 310700 700
rect 319600 500 319800 700
rect 330500 6300 330700 6500
rect 339300 6300 339500 6500
rect 340500 6300 340700 6500
rect 349600 6300 349800 6500
rect 337300 3900 337500 4300
rect 342700 3900 342900 4300
rect 339920 3640 340080 3680
rect 339920 3560 339960 3640
rect 340040 3560 340080 3640
rect 339920 3520 340080 3560
rect 337300 2900 337500 3300
rect 342700 2900 342900 3300
rect 330500 500 330700 700
rect 339300 500 339500 700
rect 340500 500 340700 700
rect 349600 500 349800 700
rect 360500 6300 360700 6500
rect 369300 6300 369500 6500
rect 370500 6300 370700 6500
rect 379600 6300 379800 6500
rect 367300 3900 367500 4300
rect 372700 3900 372900 4300
rect 369920 3640 370080 3680
rect 369920 3560 369960 3640
rect 370040 3560 370080 3640
rect 369920 3520 370080 3560
rect 367300 2900 367500 3300
rect 372700 2900 372900 3300
rect 360500 500 360700 700
rect 369300 500 369500 700
rect 370500 500 370700 700
rect 379600 500 379800 700
<< psubdiffcont >>
rect 30300 6800 50000 6900
rect 30100 300 30200 6700
rect 50100 300 50200 6700
rect 30300 100 50000 200
rect 60300 6800 80000 6900
rect 60100 300 60200 6700
rect 80100 300 80200 6700
rect 60300 100 80000 200
rect 90300 6800 110000 6900
rect 90100 300 90200 6700
rect 110100 300 110200 6700
rect 90300 100 110000 200
rect 120300 6800 140000 6900
rect 120100 300 120200 6700
rect 140100 300 140200 6700
rect 120300 100 140000 200
rect 150300 6800 170000 6900
rect 150100 300 150200 6700
rect 170100 300 170200 6700
rect 150300 100 170000 200
rect 180300 6800 200000 6900
rect 180100 300 180200 6700
rect 200100 300 200200 6700
rect 180300 100 200000 200
rect 210300 6800 230000 6900
rect 210100 300 210200 6700
rect 230100 300 230200 6700
rect 210300 100 230000 200
rect 240300 6800 260000 6900
rect 240100 300 240200 6700
rect 260100 300 260200 6700
rect 240300 100 260000 200
rect 270300 6800 290000 6900
rect 270100 300 270200 6700
rect 290100 300 290200 6700
rect 270300 100 290000 200
rect 300300 6800 320000 6900
rect 300100 300 300200 6700
rect 320100 300 320200 6700
rect 300300 100 320000 200
rect 330300 6800 350000 6900
rect 330100 300 330200 6700
rect 350100 300 350200 6700
rect 330300 100 350000 200
rect 360300 6800 380000 6900
rect 360100 300 360200 6700
rect 380100 300 380200 6700
rect 360300 100 380000 200
<< nsubdiffcont >>
rect 39500 6300 40500 6500
rect 30500 700 30700 6300
rect 37300 3300 37500 3900
rect 39960 3560 40040 3640
rect 42700 3300 42900 3900
rect 49600 700 49800 6300
rect 39500 500 40500 700
rect 69500 6300 70500 6500
rect 60500 700 60700 6300
rect 67300 3300 67500 3900
rect 69960 3560 70040 3640
rect 72700 3300 72900 3900
rect 79600 700 79800 6300
rect 69500 500 70500 700
rect 99500 6300 100500 6500
rect 90500 700 90700 6300
rect 97300 3300 97500 3900
rect 99960 3560 100040 3640
rect 102700 3300 102900 3900
rect 109600 700 109800 6300
rect 99500 500 100500 700
rect 129500 6300 130500 6500
rect 120500 700 120700 6300
rect 127300 3300 127500 3900
rect 129960 3560 130040 3640
rect 132700 3300 132900 3900
rect 139600 700 139800 6300
rect 129500 500 130500 700
rect 159500 6300 160500 6500
rect 150500 700 150700 6300
rect 157300 3300 157500 3900
rect 159960 3560 160040 3640
rect 162700 3300 162900 3900
rect 169600 700 169800 6300
rect 159500 500 160500 700
rect 189500 6300 190500 6500
rect 180500 700 180700 6300
rect 187300 3300 187500 3900
rect 189960 3560 190040 3640
rect 192700 3300 192900 3900
rect 199600 700 199800 6300
rect 189500 500 190500 700
rect 219500 6300 220500 6500
rect 210500 700 210700 6300
rect 217300 3300 217500 3900
rect 219960 3560 220040 3640
rect 222700 3300 222900 3900
rect 229600 700 229800 6300
rect 219500 500 220500 700
rect 249500 6300 250500 6500
rect 240500 700 240700 6300
rect 247300 3300 247500 3900
rect 249960 3560 250040 3640
rect 252700 3300 252900 3900
rect 259600 700 259800 6300
rect 249500 500 250500 700
rect 279500 6300 280500 6500
rect 270500 700 270700 6300
rect 277300 3300 277500 3900
rect 279960 3560 280040 3640
rect 282700 3300 282900 3900
rect 289600 700 289800 6300
rect 279500 500 280500 700
rect 309500 6300 310500 6500
rect 300500 700 300700 6300
rect 307300 3300 307500 3900
rect 309960 3560 310040 3640
rect 312700 3300 312900 3900
rect 319600 700 319800 6300
rect 309500 500 310500 700
rect 339500 6300 340500 6500
rect 330500 700 330700 6300
rect 337300 3300 337500 3900
rect 339960 3560 340040 3640
rect 342700 3300 342900 3900
rect 349600 700 349800 6300
rect 339500 500 340500 700
rect 369500 6300 370500 6500
rect 360500 700 360700 6300
rect 367300 3300 367500 3900
rect 369960 3560 370040 3640
rect 372700 3300 372900 3900
rect 379600 700 379800 6300
rect 369500 500 370500 700
<< locali >>
rect 51700 7600 52500 8700
rect 30100 6900 380500 7600
rect 30100 6800 30300 6900
rect 50000 6800 60300 6900
rect 80000 6800 90300 6900
rect 110000 6800 120300 6900
rect 140000 6800 150300 6900
rect 170000 6800 180300 6900
rect 200000 6800 210300 6900
rect 230000 6800 240300 6900
rect 260000 6800 270300 6900
rect 290000 6800 300300 6900
rect 320000 6800 330300 6900
rect 350000 6800 360300 6900
rect 380000 6800 380500 6900
rect 30100 6700 30200 6800
rect 50100 6700 50200 6800
rect 30500 6300 30700 6500
rect 39300 6300 39500 6500
rect 40500 6300 40700 6500
rect 49600 6300 49800 6500
rect 37300 3900 37500 4300
rect 42700 3900 42900 4300
rect 39900 3640 40100 3700
rect 39900 3560 39960 3640
rect 40040 3560 40100 3640
rect 39900 3500 40100 3560
rect 37300 2900 37500 3300
rect 39950 1230 40050 3500
rect 42700 2900 42900 3300
rect 39950 1130 41080 1230
rect 30500 500 30700 700
rect 39300 500 39500 700
rect 40500 500 40700 700
rect 40980 400 41080 1130
rect 49600 500 49800 700
rect 30100 200 30200 300
rect 50100 200 50200 300
rect 30100 100 30300 200
rect 50000 100 50200 200
rect 60100 6700 60200 6800
rect 80100 6700 80200 6800
rect 60500 6300 60700 6500
rect 69300 6300 69500 6500
rect 70500 6300 70700 6500
rect 79600 6300 79800 6500
rect 67300 3900 67500 4300
rect 72700 3900 72900 4300
rect 69920 3640 70080 3680
rect 69920 3560 69960 3640
rect 70040 3560 70080 3640
rect 69920 3520 70080 3560
rect 67300 2900 67500 3300
rect 69935 1765 70065 3520
rect 72700 2900 72900 3300
rect 69935 1635 70930 1765
rect 60500 500 60700 700
rect 69300 500 69500 700
rect 70500 500 70700 700
rect 70800 599 70930 1635
rect 70800 481 70806 599
rect 70924 481 70930 599
rect 79600 500 79800 700
rect 70800 475 70930 481
rect 60100 200 60200 300
rect 80100 200 80200 300
rect 60100 100 60300 200
rect 80000 100 80200 200
rect 90100 6700 90200 6800
rect 110100 6700 110200 6800
rect 90500 6300 90700 6500
rect 99300 6300 99500 6500
rect 100500 6300 100700 6500
rect 109600 6300 109800 6500
rect 97300 3900 97500 4300
rect 102700 3900 102900 4300
rect 99920 3640 100080 3680
rect 99920 3560 99960 3640
rect 100040 3560 100080 3640
rect 99920 3520 100080 3560
rect 97300 2900 97500 3300
rect 99960 830 100040 3520
rect 102700 2900 102900 3300
rect 99960 750 100810 830
rect 90500 500 90700 700
rect 99300 500 99500 700
rect 100500 500 100700 700
rect 109600 500 109800 700
rect 90100 200 90200 300
rect 110100 200 110200 300
rect 90100 100 90300 200
rect 110000 100 110200 200
rect 120100 6700 120200 6800
rect 140100 6700 140200 6800
rect 120500 6300 120700 6500
rect 129300 6300 129500 6500
rect 130500 6300 130700 6500
rect 139600 6300 139800 6500
rect 127300 3900 127500 4300
rect 132700 3900 132900 4300
rect 129920 3640 130080 3680
rect 129920 3560 129960 3640
rect 130040 3560 130080 3640
rect 129920 3520 130080 3560
rect 127300 2900 127500 3300
rect 129960 830 130040 3520
rect 132700 2900 132900 3300
rect 120500 500 120700 700
rect 129300 500 129500 700
rect 130500 500 130700 700
rect 139600 500 139800 700
rect 120100 200 120200 300
rect 140100 200 140200 300
rect 120100 100 120300 200
rect 140000 100 140200 200
rect 150100 6700 150200 6800
rect 170100 6700 170200 6800
rect 150500 6300 150700 6500
rect 159300 6300 159500 6500
rect 160500 6300 160700 6500
rect 169600 6300 169800 6500
rect 157300 3900 157500 4300
rect 162700 3900 162900 4300
rect 159920 3640 160080 3680
rect 159920 3560 159960 3640
rect 160040 3560 160080 3640
rect 159920 3520 160080 3560
rect 157300 2900 157500 3300
rect 159960 880 160040 3520
rect 162700 2900 162900 3300
rect 159960 800 161140 880
rect 150500 500 150700 700
rect 159300 500 159500 700
rect 160500 500 160700 700
rect 161060 600 161140 800
rect 169600 500 169800 700
rect 150100 200 150200 300
rect 170100 200 170200 300
rect 150100 100 150300 200
rect 170000 100 170200 200
rect 180100 6700 180200 6800
rect 200100 6700 200200 6800
rect 180500 6300 180700 6500
rect 189300 6300 189500 6500
rect 190500 6300 190700 6500
rect 199600 6300 199800 6500
rect 187300 3900 187500 4300
rect 192700 3900 192900 4300
rect 189920 3640 190080 3680
rect 189920 3560 189960 3640
rect 190040 3560 190080 3640
rect 189920 3520 190080 3560
rect 187300 2900 187500 3300
rect 189960 840 190040 3520
rect 192700 2900 192900 3300
rect 189960 760 191140 840
rect 180500 500 180700 700
rect 189300 500 189500 700
rect 190500 500 190700 700
rect 191060 580 191140 760
rect 199600 500 199800 700
rect 180100 200 180200 300
rect 200100 200 200200 300
rect 180100 100 180300 200
rect 200000 100 200200 200
rect 210100 6700 210200 6800
rect 230100 6700 230200 6800
rect 210500 6300 210700 6500
rect 219300 6300 219500 6500
rect 220500 6300 220700 6500
rect 229600 6300 229800 6500
rect 217300 3900 217500 4300
rect 222700 3900 222900 4300
rect 219920 3640 220080 3680
rect 219920 3560 219960 3640
rect 220040 3560 220080 3640
rect 219920 3520 220080 3560
rect 217300 2900 217500 3300
rect 219960 840 220040 3520
rect 222700 2900 222900 3300
rect 219960 760 221140 840
rect 210500 500 210700 700
rect 219300 500 219500 700
rect 220500 500 220700 700
rect 221060 550 221140 760
rect 229600 500 229800 700
rect 210100 200 210200 300
rect 230100 200 230200 300
rect 210100 100 210300 200
rect 230000 100 230200 200
rect 240100 6700 240200 6800
rect 260100 6700 260200 6800
rect 240500 6300 240700 6500
rect 249300 6300 249500 6500
rect 250500 6300 250700 6500
rect 259600 6300 259800 6500
rect 247300 3900 247500 4300
rect 252700 3900 252900 4300
rect 249920 3640 250080 3680
rect 249920 3560 249960 3640
rect 250040 3560 250080 3640
rect 249920 3520 250080 3560
rect 247300 2900 247500 3300
rect 249960 820 250040 3520
rect 252700 2900 252900 3300
rect 249960 740 251130 820
rect 240500 500 240700 700
rect 249300 500 249500 700
rect 250500 500 250700 700
rect 251050 480 251130 740
rect 259600 500 259800 700
rect 240100 200 240200 300
rect 260100 200 260200 300
rect 240100 100 240300 200
rect 260000 100 260200 200
rect 270100 6700 270200 6800
rect 290100 6700 290200 6800
rect 270500 6300 270700 6500
rect 279300 6300 279500 6500
rect 280500 6300 280700 6500
rect 289600 6300 289800 6500
rect 277300 3900 277500 4300
rect 282700 3900 282900 4300
rect 279920 3640 280080 3680
rect 279920 3560 279960 3640
rect 280040 3560 280080 3640
rect 279920 3520 280080 3560
rect 277300 2900 277500 3300
rect 279960 820 280040 3520
rect 282700 2900 282900 3300
rect 279960 740 281130 820
rect 270500 500 270700 700
rect 279300 500 279500 700
rect 280500 500 280700 700
rect 281050 480 281130 740
rect 289600 500 289800 700
rect 270100 200 270200 300
rect 290100 200 290200 300
rect 270100 100 270300 200
rect 290000 100 290200 200
rect 300100 6700 300200 6800
rect 320100 6700 320200 6800
rect 300500 6300 300700 6500
rect 309300 6300 309500 6500
rect 310500 6300 310700 6500
rect 319600 6300 319800 6500
rect 307300 3900 307500 4300
rect 312700 3900 312900 4300
rect 309920 3640 310080 3680
rect 309920 3560 309960 3640
rect 310040 3560 310080 3640
rect 309920 3520 310080 3560
rect 307300 2900 307500 3300
rect 309960 820 310040 3520
rect 312700 2900 312900 3300
rect 309960 740 311130 820
rect 300500 500 300700 700
rect 309300 500 309500 700
rect 310500 500 310700 700
rect 311050 480 311130 740
rect 319600 500 319800 700
rect 300100 200 300200 300
rect 320100 200 320200 300
rect 300100 100 300300 200
rect 320000 100 320200 200
rect 330100 6700 330200 6800
rect 350100 6700 350200 6800
rect 330500 6300 330700 6500
rect 339300 6300 339500 6500
rect 340500 6300 340700 6500
rect 349600 6300 349800 6500
rect 337300 3900 337500 4300
rect 342700 3900 342900 4300
rect 339920 3640 340080 3680
rect 339920 3560 339960 3640
rect 340040 3560 340080 3640
rect 339920 3520 340080 3560
rect 337300 2900 337500 3300
rect 339960 820 340040 3520
rect 342700 2900 342900 3300
rect 339960 740 341130 820
rect 330500 500 330700 700
rect 339300 500 339500 700
rect 340500 500 340700 700
rect 341050 480 341130 740
rect 349600 500 349800 700
rect 330100 200 330200 300
rect 350100 200 350200 300
rect 330100 100 330300 200
rect 350000 100 350200 200
rect 360100 6700 360200 6800
rect 380100 6700 380200 6800
rect 360500 6300 360700 6500
rect 369300 6300 369500 6500
rect 370500 6300 370700 6500
rect 379600 6300 379800 6500
rect 367300 3900 367500 4300
rect 372700 3900 372900 4300
rect 369920 3640 370080 3680
rect 369920 3560 369960 3640
rect 370040 3560 370080 3640
rect 369920 3520 370080 3560
rect 367300 2900 367500 3300
rect 369960 820 370040 3520
rect 372700 2900 372900 3300
rect 369960 740 371130 820
rect 360500 500 360700 700
rect 369300 500 369500 700
rect 370500 500 370700 700
rect 371050 480 371130 740
rect 379600 500 379800 700
rect 360100 200 360200 300
rect 380100 200 380200 300
rect 360100 100 360300 200
rect 380000 100 380200 200
<< viali >>
rect 51700 8700 52500 9500
rect 40980 300 41080 400
rect 70806 481 70924 599
rect 100810 750 100890 830
rect 129960 750 130040 830
rect 161060 520 161140 600
rect 191060 500 191140 580
rect 221060 470 221140 550
rect 251050 400 251130 480
rect 281050 400 281130 480
rect 311050 400 311130 480
rect 341050 400 341130 480
rect 371050 400 371130 480
<< metal1 >>
rect 51694 9506 52506 9512
rect 51688 8706 51694 9506
rect 52506 8706 52512 9506
rect 51688 8700 51700 8706
rect 52500 8700 52512 8706
rect 51688 8694 52512 8700
rect 100798 830 100902 836
rect 100798 750 100810 830
rect 100890 750 100902 830
rect 100798 744 100902 750
rect 129948 830 130052 836
rect 129948 750 129960 830
rect 130040 750 130890 830
rect 129948 744 130052 750
rect 70800 599 70930 611
rect 70800 481 70806 599
rect 70924 481 70930 599
rect 40968 400 41092 406
rect 40968 300 40980 400
rect 41080 300 41092 400
rect 40968 294 41092 300
rect 40980 -1150 41080 294
rect 70800 -450 70930 481
rect 100810 0 100890 744
rect 130810 0 130890 750
rect 161048 600 161152 606
rect 161048 520 161060 600
rect 161140 520 161152 600
rect 161048 514 161152 520
rect 191048 580 191152 586
rect 100800 -350 100890 0
rect 130800 -100 130890 0
rect 161060 -90 161140 514
rect 191048 500 191060 580
rect 191140 500 191152 580
rect 191048 494 191152 500
rect 221048 550 221152 556
rect 191060 -90 191140 494
rect 221048 470 221060 550
rect 221140 470 221152 550
rect 221048 464 221152 470
rect 251038 480 251142 486
rect 221060 -90 221140 464
rect 251038 400 251050 480
rect 251130 400 251142 480
rect 251038 394 251142 400
rect 281038 480 281142 486
rect 281038 400 281050 480
rect 281130 400 281142 480
rect 281038 394 281142 400
rect 311038 480 311142 486
rect 311038 400 311050 480
rect 311130 400 311142 480
rect 311038 394 311142 400
rect 341038 480 341142 486
rect 341038 400 341050 480
rect 341130 400 341142 480
rect 341038 394 341142 400
rect 371038 480 371142 486
rect 371038 400 371050 480
rect 371130 400 371142 480
rect 371038 394 371142 400
rect 251050 -90 251130 394
rect 281050 -90 281130 394
rect 311050 -90 311130 394
rect 341050 -90 341130 394
rect 371050 -90 371130 394
rect 161040 -100 161160 -90
rect 130800 -200 131150 -100
rect 161040 -120 161050 -100
rect 101050 -350 101150 -344
rect 71050 -450 71150 -444
rect 100800 -450 101050 -350
rect 70800 -550 71050 -450
rect 101050 -456 101150 -450
rect 71050 -556 71150 -550
rect 131050 -700 131150 -200
rect 161150 -120 161160 -100
rect 191040 -100 191160 -90
rect 191040 -120 191050 -100
rect 161050 -206 161150 -200
rect 191150 -120 191160 -100
rect 221040 -100 221160 -90
rect 191050 -206 191150 -200
rect 221040 -200 221050 -100
rect 221150 -200 221160 -100
rect 221040 -210 221160 -200
rect 251040 -100 251160 -90
rect 251040 -200 251050 -100
rect 251150 -200 251160 -100
rect 251040 -210 251160 -200
rect 281040 -100 281160 -90
rect 281040 -200 281050 -100
rect 281150 -200 281160 -100
rect 281040 -210 281160 -200
rect 311040 -100 311160 -90
rect 311040 -200 311050 -100
rect 311150 -200 311160 -100
rect 311040 -210 311160 -200
rect 341040 -100 341160 -90
rect 341040 -200 341050 -100
rect 341150 -200 341160 -100
rect 341040 -210 341160 -200
rect 371040 -100 371160 -90
rect 371040 -200 371050 -100
rect 371150 -200 371160 -100
rect 371040 -210 371160 -200
rect 131050 -806 131150 -800
rect 40980 -1256 41080 -1250
<< via1 >>
rect 51694 9500 52506 9506
rect 51694 8706 51700 9500
rect 51700 8706 52500 9500
rect 52500 8706 52506 9500
rect 101050 -450 101150 -350
rect 71050 -550 71150 -450
rect 161050 -200 161150 -100
rect 191050 -200 191150 -100
rect 221050 -200 221150 -100
rect 251050 -200 251150 -100
rect 281050 -200 281150 -100
rect 311050 -200 311150 -100
rect 341050 -200 341150 -100
rect 371050 -200 371150 -100
rect 131050 -800 131150 -700
rect 40980 -1250 41080 -1150
<< obsm1 >>
rect 30900 900 49400 6100
rect 60900 900 79400 6100
rect 91500 900 108800 6100
rect 121500 900 138800 6100
rect 152100 900 168200 6100
rect 182100 900 198200 6100
rect 212700 900 227600 6100
rect 242700 900 257600 6100
rect 272700 900 287600 6100
rect 302700 900 317600 6100
rect 332700 900 347600 6100
rect 362700 900 377600 6100
<< metal2 >>
rect 51600 9506 52600 9600
rect 51600 8706 51694 9506
rect 52506 8706 52600 9506
rect 51600 8600 52600 8706
rect 221050 -100 221150 -94
rect 161044 -200 161050 -100
rect 161150 -200 161156 -100
rect 191044 -200 191050 -100
rect 191150 -200 191156 -100
rect 101044 -450 101050 -350
rect 101150 -450 101156 -350
rect 71044 -550 71050 -450
rect 71150 -550 71156 -450
rect 71050 -900 71150 -550
rect 101050 -900 101150 -450
rect 131044 -800 131050 -700
rect 131150 -800 131156 -700
rect 131050 -900 131150 -800
rect 161050 -900 161150 -200
rect 191050 -900 191150 -200
rect 221050 -900 221150 -200
rect 251050 -100 251150 -94
rect 251050 -900 251150 -200
rect 281050 -100 281150 -94
rect 281050 -900 281150 -200
rect 311050 -100 311150 -94
rect 311050 -900 311150 -200
rect 341050 -100 341150 -94
rect 341050 -900 341150 -200
rect 371050 -100 371150 -94
rect 371050 -900 371150 -200
rect 71000 -1000 71200 -900
rect 101000 -1000 101200 -900
rect 131000 -1000 131200 -900
rect 161000 -1000 161200 -900
rect 191000 -1000 191200 -900
rect 221000 -1000 221200 -900
rect 251000 -1000 251200 -900
rect 281000 -1000 281200 -900
rect 311000 -1000 311200 -900
rect 341000 -1000 341200 -900
rect 371000 -1000 371200 -900
rect 40500 -1150 41750 -1000
rect 40500 -1250 40980 -1150
rect 41080 -1250 41750 -1150
rect 40500 -2000 41750 -1250
rect 70500 -2000 71750 -1000
rect 100500 -2000 101750 -1000
rect 130500 -2000 131750 -1000
rect 160500 -2000 161750 -1000
rect 190500 -2000 191750 -1000
rect 220500 -2000 221750 -1000
rect 250500 -2000 251750 -1000
rect 280500 -2000 281750 -1000
rect 310500 -2000 311750 -1000
rect 340500 -2000 341750 -1000
rect 370500 -2000 371750 -1000
<< via2 >>
rect 51694 8706 52506 9506
<< obsm2 >>
rect 30000 0 50300 7100
rect 60000 0 80400 7200
rect 90000 0 110400 7200
rect 120000 0 140400 7200
rect 150000 0 170400 7200
rect 180000 0 200400 7200
rect 210000 0 230400 7200
rect 240000 0 260400 7200
rect 270000 0 290400 7200
rect 300000 0 320400 7200
rect 330000 0 350400 7200
rect 360000 0 380400 7200
<< metal3 >>
rect 51600 9511 52600 9600
rect 51600 8701 51689 9511
rect 52511 8701 52600 9511
rect 51600 8600 52600 8701
<< obsm3 >>
rect 30000 0 50300 7100
rect 60000 0 80400 7200
rect 90000 0 110400 7200
rect 120000 0 140400 7200
rect 150000 0 170400 7200
rect 180000 0 200400 7200
rect 210000 0 230400 7200
rect 240000 0 260400 7200
rect 270000 0 290400 7200
rect 300000 0 320400 7200
rect 330000 0 350400 7200
rect 360000 0 380400 7200
<< via3 >>
rect 51689 9506 52511 9511
rect 51689 8706 51694 9506
rect 51694 8706 52506 9506
rect 52506 8706 52511 9506
rect 51689 8701 52511 8706
<< metal4 >>
rect 49300 13400 54100 14200
rect 49300 12828 54094 13400
rect 49292 12600 54094 12828
rect 49292 11890 54082 12600
rect 49282 9511 55300 9858
rect 49282 9450 51689 9511
rect 49300 8701 51689 9450
rect 52511 8701 55300 9511
rect 49300 8700 55300 8701
<< obsm4 >>
rect 30000 0 50300 7100
rect 60000 0 80400 7200
rect 90000 0 110400 7200
rect 120000 0 140400 7200
rect 150000 0 170400 7200
rect 180000 0 200400 7200
rect 210000 0 230400 7200
rect 240000 0 260400 7200
rect 270000 0 290400 7200
rect 300000 0 320400 7200
rect 330000 0 350400 7200
rect 360000 0 380400 7200
<< fillblock >>
rect 30200 200 50000 6800
rect 60200 200 80000 6800
rect 90200 200 110000 6800
rect 120200 200 140000 6800
rect 150200 200 170000 6800
rect 180200 200 200000 6800
rect 210200 200 230000 6800
rect 240200 200 260000 6800
rect 270200 200 290000 6800
rect 300200 200 320000 6800
rect 330200 200 350000 6800
rect 360200 200 380000 6800
<< labels >>
flabel metal2 41000 -1750 41000 -1750 0 FreeSans 1600 0 0 0 PD1
port 0 nsew default input
flabel metal2 71000 -1750 71000 -1750 0 FreeSans 1600 0 0 0 PD2
port 1 nsew default input
flabel metal2 101000 -1750 101000 -1750 0 FreeSans 1600 0 0 0 PD3
port 2 nsew default input
flabel metal2 131000 -1750 131000 -1750 0 FreeSans 1600 0 0 0 PD4
port 3 nsew default input
flabel metal2 161000 -1750 161000 -1750 0 FreeSans 1600 0 0 0 PD5
port 4 nsew default input
flabel metal2 191000 -1750 191000 -1750 0 FreeSans 1600 0 0 0 PD6
port 5 nsew default input
flabel metal2 221000 -1750 221000 -1750 0 FreeSans 1600 0 0 0 PD7
port 6 nsew default input
flabel metal2 251000 -1750 251000 -1750 0 FreeSans 1600 0 0 0 PD8
port 7 nsew default input
flabel metal2 281000 -1750 281000 -1750 0 FreeSans 1600 0 0 0 PD9
port 8 nsew default input
flabel metal2 311000 -1750 311000 -1750 0 FreeSans 1600 0 0 0 PD10
port 9 nsew default input
flabel metal2 341000 -1750 341000 -1750 0 FreeSans 1600 0 0 0 PD11
port 10 nsew default input
flabel metal2 371000 -1750 371000 -1750 0 FreeSans 1600 0 0 0 PD12
port 11 nsew default input
flabel metal4 49500 9250 49500 9250 0 FreeSans 1600 0 0 0 VSS
port 12 nsew ground input
flabel metal4 50900 13400 52100 14000 0 FreeSans 1600 0 0 0 VDD
port 14 nsew power input
<< end >>
